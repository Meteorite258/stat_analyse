module aes_128(clk,  state, key, out);
wire  [127:0] _000_;
input  clk;
wire  [127:0] k0;
wire  [127:0] k0b;
wire  [127:0] k1;
wire  [127:0] k1b;
wire  [127:0] k2;
wire  [127:0] k2b;
wire  [127:0] k3;
wire  [127:0] k3b;
wire  [127:0] k4;
wire  [127:0] k4b;
wire  [127:0] k5;
wire  [127:0] k5b;
wire  [127:0] k6;
wire  [127:0] k6b;
wire  [127:0] k7;
wire  [127:0] k7b;
wire  [127:0] k8;
wire  [127:0] k8b;
wire  [127:0] k9;
wire  [127:0] k9b;
input  [127:0] key;
output  [127:0] out;
wire  [127:0] s0;
wire  [127:0] s1;
wire  [127:0] s2;
wire  [127:0] s3;
wire  [127:0] s4;
wire  [127:0] s5;
wire  [127:0] s6;
wire  [127:0] s7;
wire  [127:0] s8;
wire  [127:0] s9;
input  [127:0] state;
LUT2  #(
    .INIT(4'h6)
  ) _001_ (
    .I0(state[0]),
    .I1(key[0]),
    .O(_000_[0])
  );
LUT2  #(
    .INIT(4'h6)
  ) _002_ (
    .I0(state[1]),
    .I1(key[1]),
    .O(_000_[1])
  );
LUT2  #(
    .INIT(4'h6)
  ) _003_ (
    .I0(state[2]),
    .I1(key[2]),
    .O(_000_[2])
  );
LUT2  #(
    .INIT(4'h6)
  ) _004_ (
    .I0(state[3]),
    .I1(key[3]),
    .O(_000_[3])
  );
LUT2  #(
    .INIT(4'h6)
  ) _005_ (
    .I0(state[4]),
    .I1(key[4]),
    .O(_000_[4])
  );
LUT2  #(
    .INIT(4'h6)
  ) _006_ (
    .I0(state[5]),
    .I1(key[5]),
    .O(_000_[5])
  );
LUT2  #(
    .INIT(4'h6)
  ) _007_ (
    .I0(state[6]),
    .I1(key[6]),
    .O(_000_[6])
  );
LUT2  #(
    .INIT(4'h6)
  ) _008_ (
    .I0(state[7]),
    .I1(key[7]),
    .O(_000_[7])
  );
LUT2  #(
    .INIT(4'h6)
  ) _009_ (
    .I0(state[8]),
    .I1(key[8]),
    .O(_000_[8])
  );
LUT2  #(
    .INIT(4'h6)
  ) _010_ (
    .I0(state[9]),
    .I1(key[9]),
    .O(_000_[9])
  );
LUT2  #(
    .INIT(4'h6)
  ) _011_ (
    .I0(state[10]),
    .I1(key[10]),
    .O(_000_[10])
  );
LUT2  #(
    .INIT(4'h6)
  ) _012_ (
    .I0(state[11]),
    .I1(key[11]),
    .O(_000_[11])
  );
LUT2  #(
    .INIT(4'h6)
  ) _013_ (
    .I0(state[12]),
    .I1(key[12]),
    .O(_000_[12])
  );
LUT2  #(
    .INIT(4'h6)
  ) _014_ (
    .I0(state[13]),
    .I1(key[13]),
    .O(_000_[13])
  );
LUT2  #(
    .INIT(4'h6)
  ) _015_ (
    .I0(state[14]),
    .I1(key[14]),
    .O(_000_[14])
  );
LUT2  #(
    .INIT(4'h6)
  ) _016_ (
    .I0(state[15]),
    .I1(key[15]),
    .O(_000_[15])
  );
LUT2  #(
    .INIT(4'h6)
  ) _017_ (
    .I0(state[16]),
    .I1(key[16]),
    .O(_000_[16])
  );
LUT2  #(
    .INIT(4'h6)
  ) _018_ (
    .I0(state[17]),
    .I1(key[17]),
    .O(_000_[17])
  );
LUT2  #(
    .INIT(4'h6)
  ) _019_ (
    .I0(state[18]),
    .I1(key[18]),
    .O(_000_[18])
  );
LUT2  #(
    .INIT(4'h6)
  ) _020_ (
    .I0(state[19]),
    .I1(key[19]),
    .O(_000_[19])
  );
LUT2  #(
    .INIT(4'h6)
  ) _021_ (
    .I0(state[20]),
    .I1(key[20]),
    .O(_000_[20])
  );
LUT2  #(
    .INIT(4'h6)
  ) _022_ (
    .I0(state[21]),
    .I1(key[21]),
    .O(_000_[21])
  );
LUT2  #(
    .INIT(4'h6)
  ) _023_ (
    .I0(state[22]),
    .I1(key[22]),
    .O(_000_[22])
  );
LUT2  #(
    .INIT(4'h6)
  ) _024_ (
    .I0(state[23]),
    .I1(key[23]),
    .O(_000_[23])
  );
LUT2  #(
    .INIT(4'h6)
  ) _025_ (
    .I0(state[24]),
    .I1(key[24]),
    .O(_000_[24])
  );
LUT2  #(
    .INIT(4'h6)
  ) _026_ (
    .I0(state[25]),
    .I1(key[25]),
    .O(_000_[25])
  );
LUT2  #(
    .INIT(4'h6)
  ) _027_ (
    .I0(state[26]),
    .I1(key[26]),
    .O(_000_[26])
  );
LUT2  #(
    .INIT(4'h6)
  ) _028_ (
    .I0(state[27]),
    .I1(key[27]),
    .O(_000_[27])
  );
LUT2  #(
    .INIT(4'h6)
  ) _029_ (
    .I0(state[28]),
    .I1(key[28]),
    .O(_000_[28])
  );
LUT2  #(
    .INIT(4'h6)
  ) _030_ (
    .I0(state[29]),
    .I1(key[29]),
    .O(_000_[29])
  );
LUT2  #(
    .INIT(4'h6)
  ) _031_ (
    .I0(state[30]),
    .I1(key[30]),
    .O(_000_[30])
  );
LUT2  #(
    .INIT(4'h6)
  ) _032_ (
    .I0(state[31]),
    .I1(key[31]),
    .O(_000_[31])
  );
LUT2  #(
    .INIT(4'h6)
  ) _033_ (
    .I0(state[32]),
    .I1(key[32]),
    .O(_000_[32])
  );
LUT2  #(
    .INIT(4'h6)
  ) _034_ (
    .I0(state[33]),
    .I1(key[33]),
    .O(_000_[33])
  );
LUT2  #(
    .INIT(4'h6)
  ) _035_ (
    .I0(state[34]),
    .I1(key[34]),
    .O(_000_[34])
  );
LUT2  #(
    .INIT(4'h6)
  ) _036_ (
    .I0(state[35]),
    .I1(key[35]),
    .O(_000_[35])
  );
LUT2  #(
    .INIT(4'h6)
  ) _037_ (
    .I0(state[36]),
    .I1(key[36]),
    .O(_000_[36])
  );
LUT2  #(
    .INIT(4'h6)
  ) _038_ (
    .I0(state[37]),
    .I1(key[37]),
    .O(_000_[37])
  );
LUT2  #(
    .INIT(4'h6)
  ) _039_ (
    .I0(state[38]),
    .I1(key[38]),
    .O(_000_[38])
  );
LUT2  #(
    .INIT(4'h6)
  ) _040_ (
    .I0(state[39]),
    .I1(key[39]),
    .O(_000_[39])
  );
LUT2  #(
    .INIT(4'h6)
  ) _041_ (
    .I0(state[40]),
    .I1(key[40]),
    .O(_000_[40])
  );
LUT2  #(
    .INIT(4'h6)
  ) _042_ (
    .I0(state[41]),
    .I1(key[41]),
    .O(_000_[41])
  );
LUT2  #(
    .INIT(4'h6)
  ) _043_ (
    .I0(state[42]),
    .I1(key[42]),
    .O(_000_[42])
  );
LUT2  #(
    .INIT(4'h6)
  ) _044_ (
    .I0(state[43]),
    .I1(key[43]),
    .O(_000_[43])
  );
LUT2  #(
    .INIT(4'h6)
  ) _045_ (
    .I0(state[44]),
    .I1(key[44]),
    .O(_000_[44])
  );
LUT2  #(
    .INIT(4'h6)
  ) _046_ (
    .I0(state[45]),
    .I1(key[45]),
    .O(_000_[45])
  );
LUT2  #(
    .INIT(4'h6)
  ) _047_ (
    .I0(state[46]),
    .I1(key[46]),
    .O(_000_[46])
  );
LUT2  #(
    .INIT(4'h6)
  ) _048_ (
    .I0(state[47]),
    .I1(key[47]),
    .O(_000_[47])
  );
LUT2  #(
    .INIT(4'h6)
  ) _049_ (
    .I0(state[48]),
    .I1(key[48]),
    .O(_000_[48])
  );
LUT2  #(
    .INIT(4'h6)
  ) _050_ (
    .I0(state[49]),
    .I1(key[49]),
    .O(_000_[49])
  );
LUT2  #(
    .INIT(4'h6)
  ) _051_ (
    .I0(state[50]),
    .I1(key[50]),
    .O(_000_[50])
  );
LUT2  #(
    .INIT(4'h6)
  ) _052_ (
    .I0(state[51]),
    .I1(key[51]),
    .O(_000_[51])
  );
LUT2  #(
    .INIT(4'h6)
  ) _053_ (
    .I0(state[52]),
    .I1(key[52]),
    .O(_000_[52])
  );
LUT2  #(
    .INIT(4'h6)
  ) _054_ (
    .I0(state[53]),
    .I1(key[53]),
    .O(_000_[53])
  );
LUT2  #(
    .INIT(4'h6)
  ) _055_ (
    .I0(state[54]),
    .I1(key[54]),
    .O(_000_[54])
  );
LUT2  #(
    .INIT(4'h6)
  ) _056_ (
    .I0(state[55]),
    .I1(key[55]),
    .O(_000_[55])
  );
LUT2  #(
    .INIT(4'h6)
  ) _057_ (
    .I0(state[56]),
    .I1(key[56]),
    .O(_000_[56])
  );
LUT2  #(
    .INIT(4'h6)
  ) _058_ (
    .I0(state[57]),
    .I1(key[57]),
    .O(_000_[57])
  );
LUT2  #(
    .INIT(4'h6)
  ) _059_ (
    .I0(state[58]),
    .I1(key[58]),
    .O(_000_[58])
  );
LUT2  #(
    .INIT(4'h6)
  ) _060_ (
    .I0(state[59]),
    .I1(key[59]),
    .O(_000_[59])
  );
LUT2  #(
    .INIT(4'h6)
  ) _061_ (
    .I0(state[60]),
    .I1(key[60]),
    .O(_000_[60])
  );
LUT2  #(
    .INIT(4'h6)
  ) _062_ (
    .I0(state[61]),
    .I1(key[61]),
    .O(_000_[61])
  );
LUT2  #(
    .INIT(4'h6)
  ) _063_ (
    .I0(state[62]),
    .I1(key[62]),
    .O(_000_[62])
  );
LUT2  #(
    .INIT(4'h6)
  ) _064_ (
    .I0(state[63]),
    .I1(key[63]),
    .O(_000_[63])
  );
LUT2  #(
    .INIT(4'h6)
  ) _065_ (
    .I0(state[64]),
    .I1(key[64]),
    .O(_000_[64])
  );
LUT2  #(
    .INIT(4'h6)
  ) _066_ (
    .I0(state[65]),
    .I1(key[65]),
    .O(_000_[65])
  );
LUT2  #(
    .INIT(4'h6)
  ) _067_ (
    .I0(state[66]),
    .I1(key[66]),
    .O(_000_[66])
  );
LUT2  #(
    .INIT(4'h6)
  ) _068_ (
    .I0(state[67]),
    .I1(key[67]),
    .O(_000_[67])
  );
LUT2  #(
    .INIT(4'h6)
  ) _069_ (
    .I0(state[68]),
    .I1(key[68]),
    .O(_000_[68])
  );
LUT2  #(
    .INIT(4'h6)
  ) _070_ (
    .I0(state[69]),
    .I1(key[69]),
    .O(_000_[69])
  );
LUT2  #(
    .INIT(4'h6)
  ) _071_ (
    .I0(state[70]),
    .I1(key[70]),
    .O(_000_[70])
  );
LUT2  #(
    .INIT(4'h6)
  ) _072_ (
    .I0(state[71]),
    .I1(key[71]),
    .O(_000_[71])
  );
LUT2  #(
    .INIT(4'h6)
  ) _073_ (
    .I0(state[72]),
    .I1(key[72]),
    .O(_000_[72])
  );
LUT2  #(
    .INIT(4'h6)
  ) _074_ (
    .I0(state[73]),
    .I1(key[73]),
    .O(_000_[73])
  );
LUT2  #(
    .INIT(4'h6)
  ) _075_ (
    .I0(state[74]),
    .I1(key[74]),
    .O(_000_[74])
  );
LUT2  #(
    .INIT(4'h6)
  ) _076_ (
    .I0(state[75]),
    .I1(key[75]),
    .O(_000_[75])
  );
LUT2  #(
    .INIT(4'h6)
  ) _077_ (
    .I0(state[76]),
    .I1(key[76]),
    .O(_000_[76])
  );
LUT2  #(
    .INIT(4'h6)
  ) _078_ (
    .I0(state[77]),
    .I1(key[77]),
    .O(_000_[77])
  );
LUT2  #(
    .INIT(4'h6)
  ) _079_ (
    .I0(state[78]),
    .I1(key[78]),
    .O(_000_[78])
  );
LUT2  #(
    .INIT(4'h6)
  ) _080_ (
    .I0(state[79]),
    .I1(key[79]),
    .O(_000_[79])
  );
LUT2  #(
    .INIT(4'h6)
  ) _081_ (
    .I0(state[80]),
    .I1(key[80]),
    .O(_000_[80])
  );
LUT2  #(
    .INIT(4'h6)
  ) _082_ (
    .I0(state[81]),
    .I1(key[81]),
    .O(_000_[81])
  );
LUT2  #(
    .INIT(4'h6)
  ) _083_ (
    .I0(state[82]),
    .I1(key[82]),
    .O(_000_[82])
  );
LUT2  #(
    .INIT(4'h6)
  ) _084_ (
    .I0(state[83]),
    .I1(key[83]),
    .O(_000_[83])
  );
LUT2  #(
    .INIT(4'h6)
  ) _085_ (
    .I0(state[84]),
    .I1(key[84]),
    .O(_000_[84])
  );
LUT2  #(
    .INIT(4'h6)
  ) _086_ (
    .I0(state[85]),
    .I1(key[85]),
    .O(_000_[85])
  );
LUT2  #(
    .INIT(4'h6)
  ) _087_ (
    .I0(state[86]),
    .I1(key[86]),
    .O(_000_[86])
  );
LUT2  #(
    .INIT(4'h6)
  ) _088_ (
    .I0(state[87]),
    .I1(key[87]),
    .O(_000_[87])
  );
LUT2  #(
    .INIT(4'h6)
  ) _089_ (
    .I0(state[88]),
    .I1(key[88]),
    .O(_000_[88])
  );
LUT2  #(
    .INIT(4'h6)
  ) _090_ (
    .I0(state[89]),
    .I1(key[89]),
    .O(_000_[89])
  );
LUT2  #(
    .INIT(4'h6)
  ) _091_ (
    .I0(state[90]),
    .I1(key[90]),
    .O(_000_[90])
  );
LUT2  #(
    .INIT(4'h6)
  ) _092_ (
    .I0(state[91]),
    .I1(key[91]),
    .O(_000_[91])
  );
LUT2  #(
    .INIT(4'h6)
  ) _093_ (
    .I0(state[92]),
    .I1(key[92]),
    .O(_000_[92])
  );
LUT2  #(
    .INIT(4'h6)
  ) _094_ (
    .I0(state[93]),
    .I1(key[93]),
    .O(_000_[93])
  );
LUT2  #(
    .INIT(4'h6)
  ) _095_ (
    .I0(state[94]),
    .I1(key[94]),
    .O(_000_[94])
  );
LUT2  #(
    .INIT(4'h6)
  ) _096_ (
    .I0(state[95]),
    .I1(key[95]),
    .O(_000_[95])
  );
LUT2  #(
    .INIT(4'h6)
  ) _097_ (
    .I0(state[96]),
    .I1(key[96]),
    .O(_000_[96])
  );
LUT2  #(
    .INIT(4'h6)
  ) _098_ (
    .I0(state[97]),
    .I1(key[97]),
    .O(_000_[97])
  );
LUT2  #(
    .INIT(4'h6)
  ) _099_ (
    .I0(state[98]),
    .I1(key[98]),
    .O(_000_[98])
  );
LUT2  #(
    .INIT(4'h6)
  ) _100_ (
    .I0(state[99]),
    .I1(key[99]),
    .O(_000_[99])
  );
LUT2  #(
    .INIT(4'h6)
  ) _101_ (
    .I0(state[100]),
    .I1(key[100]),
    .O(_000_[100])
  );
LUT2  #(
    .INIT(4'h6)
  ) _102_ (
    .I0(state[101]),
    .I1(key[101]),
    .O(_000_[101])
  );
LUT2  #(
    .INIT(4'h6)
  ) _103_ (
    .I0(state[102]),
    .I1(key[102]),
    .O(_000_[102])
  );
LUT2  #(
    .INIT(4'h6)
  ) _104_ (
    .I0(state[103]),
    .I1(key[103]),
    .O(_000_[103])
  );
LUT2  #(
    .INIT(4'h6)
  ) _105_ (
    .I0(state[104]),
    .I1(key[104]),
    .O(_000_[104])
  );
LUT2  #(
    .INIT(4'h6)
  ) _106_ (
    .I0(state[105]),
    .I1(key[105]),
    .O(_000_[105])
  );
LUT2  #(
    .INIT(4'h6)
  ) _107_ (
    .I0(state[106]),
    .I1(key[106]),
    .O(_000_[106])
  );
LUT2  #(
    .INIT(4'h6)
  ) _108_ (
    .I0(state[107]),
    .I1(key[107]),
    .O(_000_[107])
  );
LUT2  #(
    .INIT(4'h6)
  ) _109_ (
    .I0(state[108]),
    .I1(key[108]),
    .O(_000_[108])
  );
LUT2  #(
    .INIT(4'h6)
  ) _110_ (
    .I0(state[109]),
    .I1(key[109]),
    .O(_000_[109])
  );
LUT2  #(
    .INIT(4'h6)
  ) _111_ (
    .I0(state[110]),
    .I1(key[110]),
    .O(_000_[110])
  );
LUT2  #(
    .INIT(4'h6)
  ) _112_ (
    .I0(state[111]),
    .I1(key[111]),
    .O(_000_[111])
  );
LUT2  #(
    .INIT(4'h6)
  ) _113_ (
    .I0(state[112]),
    .I1(key[112]),
    .O(_000_[112])
  );
LUT2  #(
    .INIT(4'h6)
  ) _114_ (
    .I0(state[113]),
    .I1(key[113]),
    .O(_000_[113])
  );
LUT2  #(
    .INIT(4'h6)
  ) _115_ (
    .I0(state[114]),
    .I1(key[114]),
    .O(_000_[114])
  );
LUT2  #(
    .INIT(4'h6)
  ) _116_ (
    .I0(state[115]),
    .I1(key[115]),
    .O(_000_[115])
  );
LUT2  #(
    .INIT(4'h6)
  ) _117_ (
    .I0(state[116]),
    .I1(key[116]),
    .O(_000_[116])
  );
LUT2  #(
    .INIT(4'h6)
  ) _118_ (
    .I0(state[117]),
    .I1(key[117]),
    .O(_000_[117])
  );
LUT2  #(
    .INIT(4'h6)
  ) _119_ (
    .I0(state[118]),
    .I1(key[118]),
    .O(_000_[118])
  );
LUT2  #(
    .INIT(4'h6)
  ) _120_ (
    .I0(state[119]),
    .I1(key[119]),
    .O(_000_[119])
  );
LUT2  #(
    .INIT(4'h6)
  ) _121_ (
    .I0(state[120]),
    .I1(key[120]),
    .O(_000_[120])
  );
LUT2  #(
    .INIT(4'h6)
  ) _122_ (
    .I0(state[121]),
    .I1(key[121]),
    .O(_000_[121])
  );
LUT2  #(
    .INIT(4'h6)
  ) _123_ (
    .I0(state[122]),
    .I1(key[122]),
    .O(_000_[122])
  );
LUT2  #(
    .INIT(4'h6)
  ) _124_ (
    .I0(state[123]),
    .I1(key[123]),
    .O(_000_[123])
  );
LUT2  #(
    .INIT(4'h6)
  ) _125_ (
    .I0(state[124]),
    .I1(key[124]),
    .O(_000_[124])
  );
LUT2  #(
    .INIT(4'h6)
  ) _126_ (
    .I0(state[125]),
    .I1(key[125]),
    .O(_000_[125])
  );
LUT2  #(
    .INIT(4'h6)
  ) _127_ (
    .I0(state[126]),
    .I1(key[126]),
    .O(_000_[126])
  );
LUT2  #(
    .INIT(4'h6)
  ) _128_ (
    .I0(state[127]),
    .I1(key[127]),
    .O(_000_[127])
  );
FDRE  #(
    .INIT(1'hx)
  ) _129_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[0]),
    .Q(s0[0]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _130_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[1]),
    .Q(s0[1]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _131_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[2]),
    .Q(s0[2]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _132_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[3]),
    .Q(s0[3]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _133_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[4]),
    .Q(s0[4]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _134_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[5]),
    .Q(s0[5]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _135_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[6]),
    .Q(s0[6]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _136_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[7]),
    .Q(s0[7]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _137_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[8]),
    .Q(s0[8]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _138_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[9]),
    .Q(s0[9]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _139_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[10]),
    .Q(s0[10]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _140_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[11]),
    .Q(s0[11]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _141_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[12]),
    .Q(s0[12]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _142_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[13]),
    .Q(s0[13]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _143_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[14]),
    .Q(s0[14]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _144_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[15]),
    .Q(s0[15]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _145_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[16]),
    .Q(s0[16]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _146_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[17]),
    .Q(s0[17]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _147_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[18]),
    .Q(s0[18]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _148_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[19]),
    .Q(s0[19]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _149_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[20]),
    .Q(s0[20]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _150_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[21]),
    .Q(s0[21]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _151_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[22]),
    .Q(s0[22]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _152_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[23]),
    .Q(s0[23]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _153_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[24]),
    .Q(s0[24]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _154_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[25]),
    .Q(s0[25]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _155_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[26]),
    .Q(s0[26]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _156_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[27]),
    .Q(s0[27]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _157_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[28]),
    .Q(s0[28]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _158_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[29]),
    .Q(s0[29]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _159_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[30]),
    .Q(s0[30]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _160_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[31]),
    .Q(s0[31]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _161_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[32]),
    .Q(s0[32]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _162_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[33]),
    .Q(s0[33]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _163_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[34]),
    .Q(s0[34]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _164_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[35]),
    .Q(s0[35]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _165_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[36]),
    .Q(s0[36]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _166_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[37]),
    .Q(s0[37]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _167_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[38]),
    .Q(s0[38]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _168_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[39]),
    .Q(s0[39]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _169_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[40]),
    .Q(s0[40]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _170_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[41]),
    .Q(s0[41]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _171_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[42]),
    .Q(s0[42]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _172_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[43]),
    .Q(s0[43]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _173_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[44]),
    .Q(s0[44]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _174_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[45]),
    .Q(s0[45]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _175_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[46]),
    .Q(s0[46]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _176_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[47]),
    .Q(s0[47]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _177_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[48]),
    .Q(s0[48]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _178_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[49]),
    .Q(s0[49]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _179_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[50]),
    .Q(s0[50]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _180_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[51]),
    .Q(s0[51]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _181_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[52]),
    .Q(s0[52]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _182_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[53]),
    .Q(s0[53]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _183_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[54]),
    .Q(s0[54]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _184_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[55]),
    .Q(s0[55]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _185_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[56]),
    .Q(s0[56]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _186_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[57]),
    .Q(s0[57]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _187_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[58]),
    .Q(s0[58]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _188_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[59]),
    .Q(s0[59]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _189_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[60]),
    .Q(s0[60]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _190_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[61]),
    .Q(s0[61]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _191_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[62]),
    .Q(s0[62]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _192_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[63]),
    .Q(s0[63]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _193_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[64]),
    .Q(s0[64]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _194_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[65]),
    .Q(s0[65]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _195_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[66]),
    .Q(s0[66]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _196_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[67]),
    .Q(s0[67]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _197_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[68]),
    .Q(s0[68]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _198_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[69]),
    .Q(s0[69]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _199_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[70]),
    .Q(s0[70]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _200_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[71]),
    .Q(s0[71]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _201_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[72]),
    .Q(s0[72]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _202_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[73]),
    .Q(s0[73]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _203_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[74]),
    .Q(s0[74]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _204_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[75]),
    .Q(s0[75]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _205_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[76]),
    .Q(s0[76]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _206_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[77]),
    .Q(s0[77]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _207_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[78]),
    .Q(s0[78]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _208_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[79]),
    .Q(s0[79]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _209_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[80]),
    .Q(s0[80]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _210_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[81]),
    .Q(s0[81]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _211_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[82]),
    .Q(s0[82]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _212_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[83]),
    .Q(s0[83]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _213_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[84]),
    .Q(s0[84]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _214_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[85]),
    .Q(s0[85]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _215_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[86]),
    .Q(s0[86]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _216_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[87]),
    .Q(s0[87]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _217_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[88]),
    .Q(s0[88]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _218_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[89]),
    .Q(s0[89]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _219_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[90]),
    .Q(s0[90]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _220_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[91]),
    .Q(s0[91]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _221_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[92]),
    .Q(s0[92]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _222_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[93]),
    .Q(s0[93]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _223_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[94]),
    .Q(s0[94]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _224_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[95]),
    .Q(s0[95]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _225_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[96]),
    .Q(s0[96]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _226_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[97]),
    .Q(s0[97]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _227_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[98]),
    .Q(s0[98]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _228_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[99]),
    .Q(s0[99]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _229_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[100]),
    .Q(s0[100]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _230_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[101]),
    .Q(s0[101]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _231_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[102]),
    .Q(s0[102]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _232_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[103]),
    .Q(s0[103]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _233_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[104]),
    .Q(s0[104]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _234_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[105]),
    .Q(s0[105]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _235_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[106]),
    .Q(s0[106]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _236_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[107]),
    .Q(s0[107]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _237_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[108]),
    .Q(s0[108]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _238_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[109]),
    .Q(s0[109]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _239_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[110]),
    .Q(s0[110]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _240_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[111]),
    .Q(s0[111]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _241_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[112]),
    .Q(s0[112]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _242_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[113]),
    .Q(s0[113]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _243_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[114]),
    .Q(s0[114]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _244_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[115]),
    .Q(s0[115]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _245_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[116]),
    .Q(s0[116]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _246_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[117]),
    .Q(s0[117]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _247_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[118]),
    .Q(s0[118]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _248_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[119]),
    .Q(s0[119]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _249_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[120]),
    .Q(s0[120]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _250_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[121]),
    .Q(s0[121]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _251_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[122]),
    .Q(s0[122]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _252_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[123]),
    .Q(s0[123]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _253_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[124]),
    .Q(s0[124]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _254_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[125]),
    .Q(s0[125]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _255_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[126]),
    .Q(s0[126]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _256_ (
    .C(clk),
    .CE(1'h1),
    .D(_000_[127]),
    .Q(s0[127]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _257_ (
    .C(clk),
    .CE(1'h1),
    .D(key[0]),
    .Q(k0[0]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _258_ (
    .C(clk),
    .CE(1'h1),
    .D(key[1]),
    .Q(k0[1]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _259_ (
    .C(clk),
    .CE(1'h1),
    .D(key[2]),
    .Q(k0[2]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _260_ (
    .C(clk),
    .CE(1'h1),
    .D(key[3]),
    .Q(k0[3]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _261_ (
    .C(clk),
    .CE(1'h1),
    .D(key[4]),
    .Q(k0[4]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _262_ (
    .C(clk),
    .CE(1'h1),
    .D(key[5]),
    .Q(k0[5]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _263_ (
    .C(clk),
    .CE(1'h1),
    .D(key[6]),
    .Q(k0[6]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _264_ (
    .C(clk),
    .CE(1'h1),
    .D(key[7]),
    .Q(k0[7]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _265_ (
    .C(clk),
    .CE(1'h1),
    .D(key[8]),
    .Q(k0[8]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _266_ (
    .C(clk),
    .CE(1'h1),
    .D(key[9]),
    .Q(k0[9]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _267_ (
    .C(clk),
    .CE(1'h1),
    .D(key[10]),
    .Q(k0[10]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _268_ (
    .C(clk),
    .CE(1'h1),
    .D(key[11]),
    .Q(k0[11]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _269_ (
    .C(clk),
    .CE(1'h1),
    .D(key[12]),
    .Q(k0[12]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _270_ (
    .C(clk),
    .CE(1'h1),
    .D(key[13]),
    .Q(k0[13]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _271_ (
    .C(clk),
    .CE(1'h1),
    .D(key[14]),
    .Q(k0[14]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _272_ (
    .C(clk),
    .CE(1'h1),
    .D(key[15]),
    .Q(k0[15]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _273_ (
    .C(clk),
    .CE(1'h1),
    .D(key[16]),
    .Q(k0[16]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _274_ (
    .C(clk),
    .CE(1'h1),
    .D(key[17]),
    .Q(k0[17]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _275_ (
    .C(clk),
    .CE(1'h1),
    .D(key[18]),
    .Q(k0[18]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _276_ (
    .C(clk),
    .CE(1'h1),
    .D(key[19]),
    .Q(k0[19]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _277_ (
    .C(clk),
    .CE(1'h1),
    .D(key[20]),
    .Q(k0[20]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _278_ (
    .C(clk),
    .CE(1'h1),
    .D(key[21]),
    .Q(k0[21]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _279_ (
    .C(clk),
    .CE(1'h1),
    .D(key[22]),
    .Q(k0[22]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _280_ (
    .C(clk),
    .CE(1'h1),
    .D(key[23]),
    .Q(k0[23]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _281_ (
    .C(clk),
    .CE(1'h1),
    .D(key[24]),
    .Q(k0[24]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _282_ (
    .C(clk),
    .CE(1'h1),
    .D(key[25]),
    .Q(k0[25]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _283_ (
    .C(clk),
    .CE(1'h1),
    .D(key[26]),
    .Q(k0[26]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _284_ (
    .C(clk),
    .CE(1'h1),
    .D(key[27]),
    .Q(k0[27]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _285_ (
    .C(clk),
    .CE(1'h1),
    .D(key[28]),
    .Q(k0[28]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _286_ (
    .C(clk),
    .CE(1'h1),
    .D(key[29]),
    .Q(k0[29]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _287_ (
    .C(clk),
    .CE(1'h1),
    .D(key[30]),
    .Q(k0[30]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _288_ (
    .C(clk),
    .CE(1'h1),
    .D(key[31]),
    .Q(k0[31]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _289_ (
    .C(clk),
    .CE(1'h1),
    .D(key[32]),
    .Q(k0[32]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _290_ (
    .C(clk),
    .CE(1'h1),
    .D(key[33]),
    .Q(k0[33]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _291_ (
    .C(clk),
    .CE(1'h1),
    .D(key[34]),
    .Q(k0[34]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _292_ (
    .C(clk),
    .CE(1'h1),
    .D(key[35]),
    .Q(k0[35]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _293_ (
    .C(clk),
    .CE(1'h1),
    .D(key[36]),
    .Q(k0[36]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _294_ (
    .C(clk),
    .CE(1'h1),
    .D(key[37]),
    .Q(k0[37]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _295_ (
    .C(clk),
    .CE(1'h1),
    .D(key[38]),
    .Q(k0[38]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _296_ (
    .C(clk),
    .CE(1'h1),
    .D(key[39]),
    .Q(k0[39]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _297_ (
    .C(clk),
    .CE(1'h1),
    .D(key[40]),
    .Q(k0[40]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _298_ (
    .C(clk),
    .CE(1'h1),
    .D(key[41]),
    .Q(k0[41]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _299_ (
    .C(clk),
    .CE(1'h1),
    .D(key[42]),
    .Q(k0[42]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _300_ (
    .C(clk),
    .CE(1'h1),
    .D(key[43]),
    .Q(k0[43]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _301_ (
    .C(clk),
    .CE(1'h1),
    .D(key[44]),
    .Q(k0[44]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _302_ (
    .C(clk),
    .CE(1'h1),
    .D(key[45]),
    .Q(k0[45]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _303_ (
    .C(clk),
    .CE(1'h1),
    .D(key[46]),
    .Q(k0[46]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _304_ (
    .C(clk),
    .CE(1'h1),
    .D(key[47]),
    .Q(k0[47]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _305_ (
    .C(clk),
    .CE(1'h1),
    .D(key[48]),
    .Q(k0[48]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _306_ (
    .C(clk),
    .CE(1'h1),
    .D(key[49]),
    .Q(k0[49]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _307_ (
    .C(clk),
    .CE(1'h1),
    .D(key[50]),
    .Q(k0[50]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _308_ (
    .C(clk),
    .CE(1'h1),
    .D(key[51]),
    .Q(k0[51]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _309_ (
    .C(clk),
    .CE(1'h1),
    .D(key[52]),
    .Q(k0[52]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _310_ (
    .C(clk),
    .CE(1'h1),
    .D(key[53]),
    .Q(k0[53]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _311_ (
    .C(clk),
    .CE(1'h1),
    .D(key[54]),
    .Q(k0[54]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _312_ (
    .C(clk),
    .CE(1'h1),
    .D(key[55]),
    .Q(k0[55]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _313_ (
    .C(clk),
    .CE(1'h1),
    .D(key[56]),
    .Q(k0[56]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _314_ (
    .C(clk),
    .CE(1'h1),
    .D(key[57]),
    .Q(k0[57]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _315_ (
    .C(clk),
    .CE(1'h1),
    .D(key[58]),
    .Q(k0[58]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _316_ (
    .C(clk),
    .CE(1'h1),
    .D(key[59]),
    .Q(k0[59]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _317_ (
    .C(clk),
    .CE(1'h1),
    .D(key[60]),
    .Q(k0[60]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _318_ (
    .C(clk),
    .CE(1'h1),
    .D(key[61]),
    .Q(k0[61]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _319_ (
    .C(clk),
    .CE(1'h1),
    .D(key[62]),
    .Q(k0[62]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _320_ (
    .C(clk),
    .CE(1'h1),
    .D(key[63]),
    .Q(k0[63]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _321_ (
    .C(clk),
    .CE(1'h1),
    .D(key[64]),
    .Q(k0[64]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _322_ (
    .C(clk),
    .CE(1'h1),
    .D(key[65]),
    .Q(k0[65]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _323_ (
    .C(clk),
    .CE(1'h1),
    .D(key[66]),
    .Q(k0[66]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _324_ (
    .C(clk),
    .CE(1'h1),
    .D(key[67]),
    .Q(k0[67]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _325_ (
    .C(clk),
    .CE(1'h1),
    .D(key[68]),
    .Q(k0[68]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _326_ (
    .C(clk),
    .CE(1'h1),
    .D(key[69]),
    .Q(k0[69]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _327_ (
    .C(clk),
    .CE(1'h1),
    .D(key[70]),
    .Q(k0[70]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _328_ (
    .C(clk),
    .CE(1'h1),
    .D(key[71]),
    .Q(k0[71]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _329_ (
    .C(clk),
    .CE(1'h1),
    .D(key[72]),
    .Q(k0[72]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _330_ (
    .C(clk),
    .CE(1'h1),
    .D(key[73]),
    .Q(k0[73]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _331_ (
    .C(clk),
    .CE(1'h1),
    .D(key[74]),
    .Q(k0[74]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _332_ (
    .C(clk),
    .CE(1'h1),
    .D(key[75]),
    .Q(k0[75]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _333_ (
    .C(clk),
    .CE(1'h1),
    .D(key[76]),
    .Q(k0[76]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _334_ (
    .C(clk),
    .CE(1'h1),
    .D(key[77]),
    .Q(k0[77]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _335_ (
    .C(clk),
    .CE(1'h1),
    .D(key[78]),
    .Q(k0[78]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _336_ (
    .C(clk),
    .CE(1'h1),
    .D(key[79]),
    .Q(k0[79]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _337_ (
    .C(clk),
    .CE(1'h1),
    .D(key[80]),
    .Q(k0[80]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _338_ (
    .C(clk),
    .CE(1'h1),
    .D(key[81]),
    .Q(k0[81]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _339_ (
    .C(clk),
    .CE(1'h1),
    .D(key[82]),
    .Q(k0[82]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _340_ (
    .C(clk),
    .CE(1'h1),
    .D(key[83]),
    .Q(k0[83]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _341_ (
    .C(clk),
    .CE(1'h1),
    .D(key[84]),
    .Q(k0[84]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _342_ (
    .C(clk),
    .CE(1'h1),
    .D(key[85]),
    .Q(k0[85]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _343_ (
    .C(clk),
    .CE(1'h1),
    .D(key[86]),
    .Q(k0[86]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _344_ (
    .C(clk),
    .CE(1'h1),
    .D(key[87]),
    .Q(k0[87]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _345_ (
    .C(clk),
    .CE(1'h1),
    .D(key[88]),
    .Q(k0[88]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _346_ (
    .C(clk),
    .CE(1'h1),
    .D(key[89]),
    .Q(k0[89]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _347_ (
    .C(clk),
    .CE(1'h1),
    .D(key[90]),
    .Q(k0[90]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _348_ (
    .C(clk),
    .CE(1'h1),
    .D(key[91]),
    .Q(k0[91]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _349_ (
    .C(clk),
    .CE(1'h1),
    .D(key[92]),
    .Q(k0[92]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _350_ (
    .C(clk),
    .CE(1'h1),
    .D(key[93]),
    .Q(k0[93]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _351_ (
    .C(clk),
    .CE(1'h1),
    .D(key[94]),
    .Q(k0[94]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _352_ (
    .C(clk),
    .CE(1'h1),
    .D(key[95]),
    .Q(k0[95]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _353_ (
    .C(clk),
    .CE(1'h1),
    .D(key[96]),
    .Q(k0[96]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _354_ (
    .C(clk),
    .CE(1'h1),
    .D(key[97]),
    .Q(k0[97]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _355_ (
    .C(clk),
    .CE(1'h1),
    .D(key[98]),
    .Q(k0[98]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _356_ (
    .C(clk),
    .CE(1'h1),
    .D(key[99]),
    .Q(k0[99]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _357_ (
    .C(clk),
    .CE(1'h1),
    .D(key[100]),
    .Q(k0[100]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _358_ (
    .C(clk),
    .CE(1'h1),
    .D(key[101]),
    .Q(k0[101]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _359_ (
    .C(clk),
    .CE(1'h1),
    .D(key[102]),
    .Q(k0[102]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _360_ (
    .C(clk),
    .CE(1'h1),
    .D(key[103]),
    .Q(k0[103]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _361_ (
    .C(clk),
    .CE(1'h1),
    .D(key[104]),
    .Q(k0[104]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _362_ (
    .C(clk),
    .CE(1'h1),
    .D(key[105]),
    .Q(k0[105]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _363_ (
    .C(clk),
    .CE(1'h1),
    .D(key[106]),
    .Q(k0[106]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _364_ (
    .C(clk),
    .CE(1'h1),
    .D(key[107]),
    .Q(k0[107]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _365_ (
    .C(clk),
    .CE(1'h1),
    .D(key[108]),
    .Q(k0[108]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _366_ (
    .C(clk),
    .CE(1'h1),
    .D(key[109]),
    .Q(k0[109]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _367_ (
    .C(clk),
    .CE(1'h1),
    .D(key[110]),
    .Q(k0[110]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _368_ (
    .C(clk),
    .CE(1'h1),
    .D(key[111]),
    .Q(k0[111]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _369_ (
    .C(clk),
    .CE(1'h1),
    .D(key[112]),
    .Q(k0[112]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _370_ (
    .C(clk),
    .CE(1'h1),
    .D(key[113]),
    .Q(k0[113]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _371_ (
    .C(clk),
    .CE(1'h1),
    .D(key[114]),
    .Q(k0[114]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _372_ (
    .C(clk),
    .CE(1'h1),
    .D(key[115]),
    .Q(k0[115]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _373_ (
    .C(clk),
    .CE(1'h1),
    .D(key[116]),
    .Q(k0[116]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _374_ (
    .C(clk),
    .CE(1'h1),
    .D(key[117]),
    .Q(k0[117]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _375_ (
    .C(clk),
    .CE(1'h1),
    .D(key[118]),
    .Q(k0[118]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _376_ (
    .C(clk),
    .CE(1'h1),
    .D(key[119]),
    .Q(k0[119]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _377_ (
    .C(clk),
    .CE(1'h1),
    .D(key[120]),
    .Q(k0[120]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _378_ (
    .C(clk),
    .CE(1'h1),
    .D(key[121]),
    .Q(k0[121]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _379_ (
    .C(clk),
    .CE(1'h1),
    .D(key[122]),
    .Q(k0[122]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _380_ (
    .C(clk),
    .CE(1'h1),
    .D(key[123]),
    .Q(k0[123]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _381_ (
    .C(clk),
    .CE(1'h1),
    .D(key[124]),
    .Q(k0[124]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _382_ (
    .C(clk),
    .CE(1'h1),
    .D(key[125]),
    .Q(k0[125]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _383_ (
    .C(clk),
    .CE(1'h1),
    .D(key[126]),
    .Q(k0[126]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _384_ (
    .C(clk),
    .CE(1'h1),
    .D(key[127]),
    .Q(k0[127]),
    .R(1'h0)
  );
expand_key_128  a1 (
    .clk(clk),
    .in(k0),
    .out_1(k1),
    .out_2(k0b),
    .rcon(8'h01)
  );
expand_key_128  a10 (
    .clk(clk),
    .in(k9),
    .out_1(),
    .out_2(k9b),
    .rcon(8'h36)
  );
expand_key_128  a2 (
    .clk(clk),
    .in(k1),
    .out_1(k2),
    .out_2(k1b),
    .rcon(8'h02)
  );
expand_key_128  a3 (
    .clk(clk),
    .in(k2),
    .out_1(k3),
    .out_2(k2b),
    .rcon(8'h04)
  );
expand_key_128  a4 (
    .clk(clk),
    .in(k3),
    .out_1(k4),
    .out_2(k3b),
    .rcon(8'h08)
  );
expand_key_128  a5 (
    .clk(clk),
    .in(k4),
    .out_1(k5),
    .out_2(k4b),
    .rcon(8'h10)
  );
expand_key_128  a6 (
    .clk(clk),
    .in(k5),
    .out_1(k6),
    .out_2(k5b),
    .rcon(8'h20)
  );
expand_key_128  a7 (
    .clk(clk),
    .in(k6),
    .out_1(k7),
    .out_2(k6b),
    .rcon(8'h40)
  );
expand_key_128  a8 (
    .clk(clk),
    .in(k7),
    .out_1(k8),
    .out_2(k7b),
    .rcon(8'h80)
  );
expand_key_128  a9 (
    .clk(clk),
    .in(k8),
    .out_1(k9),
    .out_2(k8b),
    .rcon(8'h1b)
  );
one_round  r1 (
    .clk(clk),
    .key(k0b),
    .state_in(s0),
    .state_out(s1)
  );
one_round  r2 (
    .clk(clk),
    .key(k1b),
    .state_in(s1),
    .state_out(s2)
  );
one_round  r3 (
    .clk(clk),
    .key(k2b),
    .state_in(s2),
    .state_out(s3)
  );
one_round  r4 (
    .clk(clk),
    .key(k3b),
    .state_in(s3),
    .state_out(s4)
  );
one_round  r5 (
    .clk(clk),
    .key(k4b),
    .state_in(s4),
    .state_out(s5)
  );
one_round  r6 (
    .clk(clk),
    .key(k5b),
    .state_in(s5),
    .state_out(s6)
  );
one_round  r7 (
    .clk(clk),
    .key(k6b),
    .state_in(s6),
    .state_out(s7)
  );
one_round  r8 (
    .clk(clk),
    .key(k7b),
    .state_in(s7),
    .state_out(s8)
  );
one_round  r9 (
    .clk(clk),
    .key(k8b),
    .state_in(s8),
    .state_out(s9)
  );
final_round  rf (
    .clk(clk),
    .key_in(k9b),
    .state_in(s9),
    .state_out(out)
  );
endmodule
