module baud(sys_clk,  sys_rst_l, baud_clk);
wire  [23:0] _000_;
wire  _001_;
wire  _002_;
wire  _003_;
wire  _004_;
wire  _005_;
wire  _006_;
wire  [6:0] _007_;
wire  _008_;
wire  [6:0] _009_;
wire  _010_;
wire  [6:0] _011_;
wire  _012_;
wire  [6:0] _013_;
wire  _014_;
wire  [6:0] _015_;
wire  _016_;
wire  [6:0] _017_;
wire  _018_;
wire  [6:0] _019_;
wire  _020_;
wire  [6:0] _021_;
wire  _022_;
wire  [6:0] _023_;
wire  _024_;
wire  [6:0] _025_;
wire  _026_;
wire  [6:0] _027_;
wire  _028_;
wire  [6:0] _029_;
wire  _030_;
wire  [6:0] _031_;
wire  _032_;
wire  [6:0] _033_;
wire  _034_;
wire  [6:0] _035_;
wire  _036_;
wire  [6:0] _037_;
wire  _038_;
wire  [6:0] _039_;
wire  _040_;
wire  [6:0] _041_;
wire  _042_;
wire  [6:0] _043_;
wire  _044_;
wire  [6:0] _045_;
wire  _046_;
wire  [6:0] _047_;
wire  _048_;
wire  [6:0] _049_;
wire  _050_;
wire  [6:0] _051_;
wire  _052_;
wire  [6:0] _053_;
wire  _054_;
wire  _055_;
wire  _056_;
wire  _057_;
wire  _058_;
wire  _059_;
wire  _060_;
wire  _061_;
wire  _062_;
wire  _063_;
wire  _064_;
wire  _065_;
wire  _066_;
wire  _067_;
wire  _068_;
wire  _069_;
wire  _070_;
wire  _071_;
wire  _072_;
wire  _073_;
wire  _074_;
wire  _075_;
wire  _076_;
wire  _077_;
wire  _078_;
wire  _079_;
wire  _080_;
wire  _081_;
wire  [23:0] _082_;
wire  [23:0] _083_;
output  baud_clk;
wire  baud_clk;
wire  [23:0] clk_div;
input  sys_clk;
wire  sys_clk;
input  sys_rst_l;
wire  sys_rst_l;
LUT6  #(
    .INIT(64'h8000000000000000)
  ) _084_ (
    .I0(_007_[5]),
    .I1(_007_[0]),
    .I2(_007_[1]),
    .I3(_007_[2]),
    .I4(_007_[3]),
    .I5(_007_[4]),
    .O(_055_)
  );
MUXF7  _085_ (
    .I0(1'h0),
    .I1(1'h0),
    .O(_001_),
    .S(clk_div[10])
  );
LUT6  #(
    .INIT(64'h0000000000000001)
  ) _086_ (
    .I0(clk_div[1]),
    .I1(clk_div[3]),
    .I2(clk_div[4]),
    .I3(clk_div[5]),
    .I4(clk_div[7]),
    .I5(clk_div[9]),
    .O(_003_)
  );
MUXF7  _087_ (
    .I0(_003_),
    .I1(1'h0),
    .O(_002_),
    .S(clk_div[10])
  );
MUXF8  _088_ (
    .I0(_001_),
    .I1(_002_),
    .O(_007_[5]),
    .S(clk_div[8])
  );
LUT6  #(
    .INIT(64'h0000000000000001)
  ) _089_ (
    .I0(clk_div[11]),
    .I1(clk_div[12]),
    .I2(clk_div[13]),
    .I3(clk_div[14]),
    .I4(clk_div[15]),
    .I5(clk_div[16]),
    .O(_006_)
  );
MUXF7  _090_ (
    .I0(_006_),
    .I1(1'h0),
    .O(_004_),
    .S(clk_div[17])
  );
MUXF7  _091_ (
    .I0(1'h0),
    .I1(1'h0),
    .O(_005_),
    .S(clk_div[17])
  );
MUXF8  _092_ (
    .I0(_004_),
    .I1(_005_),
    .O(_007_[0]),
    .S(clk_div[18])
  );
LUT2  #(
    .INIT(4'h4)
  ) _093_ (
    .I0(clk_div[23]),
    .I1(clk_div[0]),
    .O(_007_[1])
  );
LUT2  #(
    .INIT(4'h8)
  ) _094_ (
    .I0(clk_div[2]),
    .I1(clk_div[6]),
    .O(_007_[2])
  );
LUT2  #(
    .INIT(4'h1)
  ) _095_ (
    .I0(clk_div[19]),
    .I1(clk_div[20]),
    .O(_007_[3])
  );
LUT2  #(
    .INIT(4'h1)
  ) _096_ (
    .I0(clk_div[21]),
    .I1(clk_div[22]),
    .O(_007_[4])
  );
LUT6  #(
    .INIT(64'h7fffffffffffffff)
  ) _097_ (
    .I0(_007_[0]),
    .I1(_007_[1]),
    .I2(_007_[2]),
    .I3(_007_[3]),
    .I4(_007_[4]),
    .I5(_007_[5]),
    .O(_008_)
  );
MUXF7  _098_ (
    .I0(1'h0),
    .I1(_008_),
    .O(_000_[0]),
    .S(_007_[6])
  );
LUT6  #(
    .INIT(64'h7fffffffffffffff)
  ) _099_ (
    .I0(_007_[0]),
    .I1(_007_[1]),
    .I2(_007_[2]),
    .I3(_007_[3]),
    .I4(_007_[4]),
    .I5(_007_[5]),
    .O(_010_)
  );
MUXF7  _100_ (
    .I0(1'h0),
    .I1(_010_),
    .O(_000_[1]),
    .S(_009_[6])
  );
LUT6  #(
    .INIT(64'h7fffffffffffffff)
  ) _101_ (
    .I0(_007_[0]),
    .I1(_007_[1]),
    .I2(_007_[2]),
    .I3(_007_[3]),
    .I4(_007_[4]),
    .I5(_007_[5]),
    .O(_012_)
  );
MUXF7  _102_ (
    .I0(1'h0),
    .I1(_012_),
    .O(_000_[2]),
    .S(_011_[6])
  );
LUT6  #(
    .INIT(64'h7fffffffffffffff)
  ) _103_ (
    .I0(_007_[0]),
    .I1(_007_[1]),
    .I2(_007_[2]),
    .I3(_007_[3]),
    .I4(_007_[4]),
    .I5(_007_[5]),
    .O(_014_)
  );
MUXF7  _104_ (
    .I0(1'h0),
    .I1(_014_),
    .O(_000_[3]),
    .S(_013_[6])
  );
LUT6  #(
    .INIT(64'h7fffffffffffffff)
  ) _105_ (
    .I0(_007_[0]),
    .I1(_007_[1]),
    .I2(_007_[2]),
    .I3(_007_[3]),
    .I4(_007_[4]),
    .I5(_007_[5]),
    .O(_016_)
  );
MUXF7  _106_ (
    .I0(1'h0),
    .I1(_016_),
    .O(_000_[4]),
    .S(_015_[6])
  );
LUT6  #(
    .INIT(64'h7fffffffffffffff)
  ) _107_ (
    .I0(_007_[0]),
    .I1(_007_[1]),
    .I2(_007_[2]),
    .I3(_007_[3]),
    .I4(_007_[4]),
    .I5(_007_[5]),
    .O(_018_)
  );
MUXF7  _108_ (
    .I0(1'h0),
    .I1(_018_),
    .O(_000_[5]),
    .S(_017_[6])
  );
LUT6  #(
    .INIT(64'h7fffffffffffffff)
  ) _109_ (
    .I0(_007_[0]),
    .I1(_007_[1]),
    .I2(_007_[2]),
    .I3(_007_[3]),
    .I4(_007_[4]),
    .I5(_007_[5]),
    .O(_020_)
  );
MUXF7  _110_ (
    .I0(1'h0),
    .I1(_020_),
    .O(_000_[6]),
    .S(_019_[6])
  );
LUT6  #(
    .INIT(64'h7fffffffffffffff)
  ) _111_ (
    .I0(_007_[0]),
    .I1(_007_[1]),
    .I2(_007_[2]),
    .I3(_007_[3]),
    .I4(_007_[4]),
    .I5(_007_[5]),
    .O(_022_)
  );
MUXF7  _112_ (
    .I0(1'h0),
    .I1(_022_),
    .O(_000_[7]),
    .S(_021_[6])
  );
LUT6  #(
    .INIT(64'h7fffffffffffffff)
  ) _113_ (
    .I0(_007_[0]),
    .I1(_007_[1]),
    .I2(_007_[2]),
    .I3(_007_[3]),
    .I4(_007_[4]),
    .I5(_007_[5]),
    .O(_024_)
  );
MUXF7  _114_ (
    .I0(1'h0),
    .I1(_024_),
    .O(_000_[8]),
    .S(_023_[6])
  );
LUT6  #(
    .INIT(64'h7fffffffffffffff)
  ) _115_ (
    .I0(_007_[0]),
    .I1(_007_[1]),
    .I2(_007_[2]),
    .I3(_007_[3]),
    .I4(_007_[4]),
    .I5(_007_[5]),
    .O(_026_)
  );
MUXF7  _116_ (
    .I0(1'h0),
    .I1(_026_),
    .O(_000_[9]),
    .S(_025_[6])
  );
LUT6  #(
    .INIT(64'h7fffffffffffffff)
  ) _117_ (
    .I0(_007_[0]),
    .I1(_007_[1]),
    .I2(_007_[2]),
    .I3(_007_[3]),
    .I4(_007_[4]),
    .I5(_007_[5]),
    .O(_028_)
  );
MUXF7  _118_ (
    .I0(1'h0),
    .I1(_028_),
    .O(_000_[10]),
    .S(_027_[6])
  );
LUT6  #(
    .INIT(64'h7fffffffffffffff)
  ) _119_ (
    .I0(_007_[0]),
    .I1(_007_[1]),
    .I2(_007_[2]),
    .I3(_007_[3]),
    .I4(_007_[4]),
    .I5(_007_[5]),
    .O(_030_)
  );
MUXF7  _120_ (
    .I0(1'h0),
    .I1(_030_),
    .O(_000_[11]),
    .S(_029_[6])
  );
LUT6  #(
    .INIT(64'h7fffffffffffffff)
  ) _121_ (
    .I0(_007_[0]),
    .I1(_007_[1]),
    .I2(_007_[2]),
    .I3(_007_[3]),
    .I4(_007_[4]),
    .I5(_007_[5]),
    .O(_032_)
  );
MUXF7  _122_ (
    .I0(1'h0),
    .I1(_032_),
    .O(_000_[12]),
    .S(_031_[6])
  );
LUT6  #(
    .INIT(64'h7fffffffffffffff)
  ) _123_ (
    .I0(_007_[0]),
    .I1(_007_[1]),
    .I2(_007_[2]),
    .I3(_007_[3]),
    .I4(_007_[4]),
    .I5(_007_[5]),
    .O(_034_)
  );
MUXF7  _124_ (
    .I0(1'h0),
    .I1(_034_),
    .O(_000_[13]),
    .S(_033_[6])
  );
LUT6  #(
    .INIT(64'h7fffffffffffffff)
  ) _125_ (
    .I0(_007_[0]),
    .I1(_007_[1]),
    .I2(_007_[2]),
    .I3(_007_[3]),
    .I4(_007_[4]),
    .I5(_007_[5]),
    .O(_036_)
  );
MUXF7  _126_ (
    .I0(1'h0),
    .I1(_036_),
    .O(_000_[14]),
    .S(_035_[6])
  );
LUT6  #(
    .INIT(64'h7fffffffffffffff)
  ) _127_ (
    .I0(_007_[0]),
    .I1(_007_[1]),
    .I2(_007_[2]),
    .I3(_007_[3]),
    .I4(_007_[4]),
    .I5(_007_[5]),
    .O(_038_)
  );
MUXF7  _128_ (
    .I0(1'h0),
    .I1(_038_),
    .O(_000_[15]),
    .S(_037_[6])
  );
LUT6  #(
    .INIT(64'h7fffffffffffffff)
  ) _129_ (
    .I0(_007_[0]),
    .I1(_007_[1]),
    .I2(_007_[2]),
    .I3(_007_[3]),
    .I4(_007_[4]),
    .I5(_007_[5]),
    .O(_040_)
  );
MUXF7  _130_ (
    .I0(1'h0),
    .I1(_040_),
    .O(_000_[16]),
    .S(_039_[6])
  );
LUT6  #(
    .INIT(64'h7fffffffffffffff)
  ) _131_ (
    .I0(_007_[0]),
    .I1(_007_[1]),
    .I2(_007_[2]),
    .I3(_007_[3]),
    .I4(_007_[4]),
    .I5(_007_[5]),
    .O(_042_)
  );
MUXF7  _132_ (
    .I0(1'h0),
    .I1(_042_),
    .O(_000_[17]),
    .S(_041_[6])
  );
LUT6  #(
    .INIT(64'h7fffffffffffffff)
  ) _133_ (
    .I0(_007_[0]),
    .I1(_007_[1]),
    .I2(_007_[2]),
    .I3(_007_[3]),
    .I4(_007_[4]),
    .I5(_007_[5]),
    .O(_044_)
  );
MUXF7  _134_ (
    .I0(1'h0),
    .I1(_044_),
    .O(_000_[18]),
    .S(_043_[6])
  );
LUT6  #(
    .INIT(64'h7fffffffffffffff)
  ) _135_ (
    .I0(_007_[0]),
    .I1(_007_[1]),
    .I2(_007_[2]),
    .I3(_007_[3]),
    .I4(_007_[4]),
    .I5(_007_[5]),
    .O(_046_)
  );
MUXF7  _136_ (
    .I0(1'h0),
    .I1(_046_),
    .O(_000_[19]),
    .S(_045_[6])
  );
LUT6  #(
    .INIT(64'h7fffffffffffffff)
  ) _137_ (
    .I0(_007_[0]),
    .I1(_007_[1]),
    .I2(_007_[2]),
    .I3(_007_[3]),
    .I4(_007_[4]),
    .I5(_007_[5]),
    .O(_048_)
  );
MUXF7  _138_ (
    .I0(1'h0),
    .I1(_048_),
    .O(_000_[20]),
    .S(_047_[6])
  );
LUT6  #(
    .INIT(64'h7fffffffffffffff)
  ) _139_ (
    .I0(_007_[0]),
    .I1(_007_[1]),
    .I2(_007_[2]),
    .I3(_007_[3]),
    .I4(_007_[4]),
    .I5(_007_[5]),
    .O(_050_)
  );
MUXF7  _140_ (
    .I0(1'h0),
    .I1(_050_),
    .O(_000_[21]),
    .S(_049_[6])
  );
LUT6  #(
    .INIT(64'h7fffffffffffffff)
  ) _141_ (
    .I0(_007_[0]),
    .I1(_007_[1]),
    .I2(_007_[2]),
    .I3(_007_[3]),
    .I4(_007_[4]),
    .I5(_007_[5]),
    .O(_052_)
  );
MUXF7  _142_ (
    .I0(1'h0),
    .I1(_052_),
    .O(_000_[22]),
    .S(_051_[6])
  );
LUT6  #(
    .INIT(64'h7fffffffffffffff)
  ) _143_ (
    .I0(_007_[0]),
    .I1(_007_[1]),
    .I2(_007_[2]),
    .I3(_007_[3]),
    .I4(_007_[4]),
    .I5(_007_[5]),
    .O(_054_)
  );
MUXF7  _144_ (
    .I0(1'h0),
    .I1(_054_),
    .O(_000_[23]),
    .S(_053_[6])
  );
INV  _145_ (
    .I(sys_rst_l),
    .O(_056_)
  );
INV  _146_ (
    .I(clk_div[0]),
    .O(_083_[0])
  );
INV  _147_ (
    .I(baud_clk),
    .O(_081_)
  );
INV  _148_ (
    .I(sys_rst_l),
    .O(_057_)
  );
INV  _149_ (
    .I(sys_rst_l),
    .O(_058_)
  );
INV  _150_ (
    .I(sys_rst_l),
    .O(_059_)
  );
INV  _151_ (
    .I(sys_rst_l),
    .O(_060_)
  );
INV  _152_ (
    .I(sys_rst_l),
    .O(_061_)
  );
INV  _153_ (
    .I(sys_rst_l),
    .O(_062_)
  );
INV  _154_ (
    .I(sys_rst_l),
    .O(_063_)
  );
INV  _155_ (
    .I(sys_rst_l),
    .O(_064_)
  );
INV  _156_ (
    .I(sys_rst_l),
    .O(_065_)
  );
INV  _157_ (
    .I(sys_rst_l),
    .O(_066_)
  );
INV  _158_ (
    .I(sys_rst_l),
    .O(_067_)
  );
INV  _159_ (
    .I(sys_rst_l),
    .O(_068_)
  );
INV  _160_ (
    .I(sys_rst_l),
    .O(_069_)
  );
INV  _161_ (
    .I(sys_rst_l),
    .O(_070_)
  );
INV  _162_ (
    .I(sys_rst_l),
    .O(_071_)
  );
INV  _163_ (
    .I(sys_rst_l),
    .O(_072_)
  );
INV  _164_ (
    .I(sys_rst_l),
    .O(_073_)
  );
INV  _165_ (
    .I(sys_rst_l),
    .O(_074_)
  );
INV  _166_ (
    .I(sys_rst_l),
    .O(_075_)
  );
INV  _167_ (
    .I(sys_rst_l),
    .O(_076_)
  );
INV  _168_ (
    .I(sys_rst_l),
    .O(_077_)
  );
INV  _169_ (
    .I(sys_rst_l),
    .O(_078_)
  );
INV  _170_ (
    .I(sys_rst_l),
    .O(_079_)
  );
INV  _171_ (
    .I(sys_rst_l),
    .O(_080_)
  );
CARRY4  _172_ (
    .CI(1'h0),
    .CO(_082_[3:0]),
    .CYINIT(1'h0),
    .DI(4'h1),
    .O({ _013_[6], _011_[6], _009_[6], _007_[6] }),
    .S({ clk_div[3:1], _083_[0] })
  );
CARRY4  _173_ (
    .CI(_082_[3]),
    .CO(_082_[7:4]),
    .CYINIT(1'h0),
    .DI(4'h0),
    .O({ _021_[6], _019_[6], _017_[6], _015_[6] }),
    .S(clk_div[7:4])
  );
CARRY4  _174_ (
    .CI(_082_[7]),
    .CO(_082_[11:8]),
    .CYINIT(1'h0),
    .DI(4'h0),
    .O({ _029_[6], _027_[6], _025_[6], _023_[6] }),
    .S(clk_div[11:8])
  );
CARRY4  _175_ (
    .CI(_082_[11]),
    .CO(_082_[15:12]),
    .CYINIT(1'h0),
    .DI(4'h0),
    .O({ _037_[6], _035_[6], _033_[6], _031_[6] }),
    .S(clk_div[15:12])
  );
CARRY4  _176_ (
    .CI(_082_[15]),
    .CO(_082_[19:16]),
    .CYINIT(1'h0),
    .DI(4'h0),
    .O({ _045_[6], _043_[6], _041_[6], _039_[6] }),
    .S(clk_div[19:16])
  );
CARRY4  _177_ (
    .CI(_082_[19]),
    .CO(_082_[23:20]),
    .CYINIT(1'h0),
    .DI(4'h0),
    .O({ _053_[6], _051_[6], _049_[6], _047_[6] }),
    .S(clk_div[23:20])
  );
FDCE  #(
    .INIT(1'hx)
  ) _178_ (
    .C(sys_clk),
    .CE(_055_),
    .CLR(_056_),
    .D(_081_),
    .Q(baud_clk)
  );
FDCE  #(
    .INIT(1'hx)
  ) _179_ (
    .C(sys_clk),
    .CE(1'h1),
    .CLR(_057_),
    .D(_000_[0]),
    .Q(clk_div[0])
  );
FDCE  #(
    .INIT(1'hx)
  ) _180_ (
    .C(sys_clk),
    .CE(1'h1),
    .CLR(_058_),
    .D(_000_[1]),
    .Q(clk_div[1])
  );
FDCE  #(
    .INIT(1'hx)
  ) _181_ (
    .C(sys_clk),
    .CE(1'h1),
    .CLR(_059_),
    .D(_000_[2]),
    .Q(clk_div[2])
  );
FDCE  #(
    .INIT(1'hx)
  ) _182_ (
    .C(sys_clk),
    .CE(1'h1),
    .CLR(_060_),
    .D(_000_[3]),
    .Q(clk_div[3])
  );
FDCE  #(
    .INIT(1'hx)
  ) _183_ (
    .C(sys_clk),
    .CE(1'h1),
    .CLR(_061_),
    .D(_000_[4]),
    .Q(clk_div[4])
  );
FDCE  #(
    .INIT(1'hx)
  ) _184_ (
    .C(sys_clk),
    .CE(1'h1),
    .CLR(_062_),
    .D(_000_[5]),
    .Q(clk_div[5])
  );
FDCE  #(
    .INIT(1'hx)
  ) _185_ (
    .C(sys_clk),
    .CE(1'h1),
    .CLR(_063_),
    .D(_000_[6]),
    .Q(clk_div[6])
  );
FDCE  #(
    .INIT(1'hx)
  ) _186_ (
    .C(sys_clk),
    .CE(1'h1),
    .CLR(_064_),
    .D(_000_[7]),
    .Q(clk_div[7])
  );
FDCE  #(
    .INIT(1'hx)
  ) _187_ (
    .C(sys_clk),
    .CE(1'h1),
    .CLR(_065_),
    .D(_000_[8]),
    .Q(clk_div[8])
  );
FDCE  #(
    .INIT(1'hx)
  ) _188_ (
    .C(sys_clk),
    .CE(1'h1),
    .CLR(_066_),
    .D(_000_[9]),
    .Q(clk_div[9])
  );
FDCE  #(
    .INIT(1'hx)
  ) _189_ (
    .C(sys_clk),
    .CE(1'h1),
    .CLR(_067_),
    .D(_000_[10]),
    .Q(clk_div[10])
  );
FDCE  #(
    .INIT(1'hx)
  ) _190_ (
    .C(sys_clk),
    .CE(1'h1),
    .CLR(_068_),
    .D(_000_[11]),
    .Q(clk_div[11])
  );
FDCE  #(
    .INIT(1'hx)
  ) _191_ (
    .C(sys_clk),
    .CE(1'h1),
    .CLR(_069_),
    .D(_000_[12]),
    .Q(clk_div[12])
  );
FDCE  #(
    .INIT(1'hx)
  ) _192_ (
    .C(sys_clk),
    .CE(1'h1),
    .CLR(_070_),
    .D(_000_[13]),
    .Q(clk_div[13])
  );
FDCE  #(
    .INIT(1'hx)
  ) _193_ (
    .C(sys_clk),
    .CE(1'h1),
    .CLR(_071_),
    .D(_000_[14]),
    .Q(clk_div[14])
  );
FDCE  #(
    .INIT(1'hx)
  ) _194_ (
    .C(sys_clk),
    .CE(1'h1),
    .CLR(_072_),
    .D(_000_[15]),
    .Q(clk_div[15])
  );
FDCE  #(
    .INIT(1'hx)
  ) _195_ (
    .C(sys_clk),
    .CE(1'h1),
    .CLR(_073_),
    .D(_000_[16]),
    .Q(clk_div[16])
  );
FDCE  #(
    .INIT(1'hx)
  ) _196_ (
    .C(sys_clk),
    .CE(1'h1),
    .CLR(_074_),
    .D(_000_[17]),
    .Q(clk_div[17])
  );
FDCE  #(
    .INIT(1'hx)
  ) _197_ (
    .C(sys_clk),
    .CE(1'h1),
    .CLR(_075_),
    .D(_000_[18]),
    .Q(clk_div[18])
  );
FDCE  #(
    .INIT(1'hx)
  ) _198_ (
    .C(sys_clk),
    .CE(1'h1),
    .CLR(_076_),
    .D(_000_[19]),
    .Q(clk_div[19])
  );
FDCE  #(
    .INIT(1'hx)
  ) _199_ (
    .C(sys_clk),
    .CE(1'h1),
    .CLR(_077_),
    .D(_000_[20]),
    .Q(clk_div[20])
  );
FDCE  #(
    .INIT(1'hx)
  ) _200_ (
    .C(sys_clk),
    .CE(1'h1),
    .CLR(_078_),
    .D(_000_[21]),
    .Q(clk_div[21])
  );
FDCE  #(
    .INIT(1'hx)
  ) _201_ (
    .C(sys_clk),
    .CE(1'h1),
    .CLR(_079_),
    .D(_000_[22]),
    .Q(clk_div[22])
  );
FDCE  #(
    .INIT(1'hx)
  ) _202_ (
    .C(sys_clk),
    .CE(1'h1),
    .CLR(_080_),
    .D(_000_[23]),
    .Q(clk_div[23])
  );
assign  _041_[5:0] = _007_[5:0];
assign  _031_[5:0] = _007_[5:0];
assign  _019_[5:0] = _007_[5:0];
assign  _023_[5:0] = _007_[5:0];
assign  _027_[5:0] = _007_[5:0];
assign  _015_[5:0] = _007_[5:0];
assign  _029_[5:0] = _007_[5:0];
assign  _039_[5:0] = _007_[5:0];
assign  _045_[5:0] = _007_[5:0];
assign  _049_[5:0] = _007_[5:0];
assign  _013_[5:0] = _007_[5:0];
assign  _037_[5:0] = _007_[5:0];
assign  _011_[5:0] = _007_[5:0];
assign  _035_[5:0] = _007_[5:0];
assign  _009_[5:0] = _007_[5:0];
assign  _043_[5:0] = _007_[5:0];
assign  _033_[5:0] = _007_[5:0];
assign  _053_[5:0] = _007_[5:0];
assign  _047_[5:0] = _007_[5:0];
assign  _025_[5:0] = _007_[5:0];
assign  _051_[5:0] = _007_[5:0];
assign  _021_[5:0] = _007_[5:0];
assign  _083_[23:1] = clk_div[23:1];
assign  _017_[5:0] = _007_[5:0];
endmodule
