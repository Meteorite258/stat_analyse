module expand_key_128(clk,  in, out_1, out_2, rcon);
input  clk;
input  [127:0] in;
wire  [31:0] k0;
wire  [31:0] k0a;
wire  [31:0] k0b;
wire  [31:0] k1;
wire  [31:0] k1a;
wire  [31:0] k1b;
wire  [31:0] k2;
wire  [31:0] k2a;
wire  [31:0] k2b;
wire  [31:0] k3;
wire  [31:0] k3a;
wire  [31:0] k3b;
wire  [31:0] k4a;
output  [127:0] out_1;
output  [127:0] out_2;
input  [7:0] rcon;
wire  [31:0] v0;
wire  [31:0] v1;
wire  [31:0] v2;
wire  [31:0] v3;
LUT2  #(
    .INIT(4'h6)
  ) _000_ (
    .I0(in[120]),
    .I1(rcon[0]),
    .O(v0[24])
  );
LUT2  #(
    .INIT(4'h6)
  ) _001_ (
    .I0(in[121]),
    .I1(rcon[1]),
    .O(v0[25])
  );
LUT2  #(
    .INIT(4'h6)
  ) _002_ (
    .I0(in[122]),
    .I1(rcon[2]),
    .O(v0[26])
  );
LUT2  #(
    .INIT(4'h6)
  ) _003_ (
    .I0(in[123]),
    .I1(rcon[3]),
    .O(v0[27])
  );
LUT2  #(
    .INIT(4'h6)
  ) _004_ (
    .I0(in[124]),
    .I1(rcon[4]),
    .O(v0[28])
  );
LUT2  #(
    .INIT(4'h6)
  ) _005_ (
    .I0(in[125]),
    .I1(rcon[5]),
    .O(v0[29])
  );
LUT2  #(
    .INIT(4'h6)
  ) _006_ (
    .I0(in[126]),
    .I1(rcon[6]),
    .O(v0[30])
  );
LUT2  #(
    .INIT(4'h6)
  ) _007_ (
    .I0(in[127]),
    .I1(rcon[7]),
    .O(v0[31])
  );
LUT2  #(
    .INIT(4'h6)
  ) _008_ (
    .I0(in[96]),
    .I1(in[64]),
    .O(v1[0])
  );
LUT2  #(
    .INIT(4'h6)
  ) _009_ (
    .I0(in[97]),
    .I1(in[65]),
    .O(v1[1])
  );
LUT2  #(
    .INIT(4'h6)
  ) _010_ (
    .I0(in[98]),
    .I1(in[66]),
    .O(v1[2])
  );
LUT2  #(
    .INIT(4'h6)
  ) _011_ (
    .I0(in[99]),
    .I1(in[67]),
    .O(v1[3])
  );
LUT2  #(
    .INIT(4'h6)
  ) _012_ (
    .I0(in[100]),
    .I1(in[68]),
    .O(v1[4])
  );
LUT2  #(
    .INIT(4'h6)
  ) _013_ (
    .I0(in[101]),
    .I1(in[69]),
    .O(v1[5])
  );
LUT2  #(
    .INIT(4'h6)
  ) _014_ (
    .I0(in[102]),
    .I1(in[70]),
    .O(v1[6])
  );
LUT2  #(
    .INIT(4'h6)
  ) _015_ (
    .I0(in[103]),
    .I1(in[71]),
    .O(v1[7])
  );
LUT2  #(
    .INIT(4'h6)
  ) _016_ (
    .I0(in[104]),
    .I1(in[72]),
    .O(v1[8])
  );
LUT2  #(
    .INIT(4'h6)
  ) _017_ (
    .I0(in[105]),
    .I1(in[73]),
    .O(v1[9])
  );
LUT2  #(
    .INIT(4'h6)
  ) _018_ (
    .I0(in[106]),
    .I1(in[74]),
    .O(v1[10])
  );
LUT2  #(
    .INIT(4'h6)
  ) _019_ (
    .I0(in[107]),
    .I1(in[75]),
    .O(v1[11])
  );
LUT2  #(
    .INIT(4'h6)
  ) _020_ (
    .I0(in[108]),
    .I1(in[76]),
    .O(v1[12])
  );
LUT2  #(
    .INIT(4'h6)
  ) _021_ (
    .I0(in[109]),
    .I1(in[77]),
    .O(v1[13])
  );
LUT2  #(
    .INIT(4'h6)
  ) _022_ (
    .I0(in[110]),
    .I1(in[78]),
    .O(v1[14])
  );
LUT2  #(
    .INIT(4'h6)
  ) _023_ (
    .I0(in[111]),
    .I1(in[79]),
    .O(v1[15])
  );
LUT2  #(
    .INIT(4'h6)
  ) _024_ (
    .I0(in[112]),
    .I1(in[80]),
    .O(v1[16])
  );
LUT2  #(
    .INIT(4'h6)
  ) _025_ (
    .I0(in[113]),
    .I1(in[81]),
    .O(v1[17])
  );
LUT2  #(
    .INIT(4'h6)
  ) _026_ (
    .I0(in[114]),
    .I1(in[82]),
    .O(v1[18])
  );
LUT2  #(
    .INIT(4'h6)
  ) _027_ (
    .I0(in[115]),
    .I1(in[83]),
    .O(v1[19])
  );
LUT2  #(
    .INIT(4'h6)
  ) _028_ (
    .I0(in[116]),
    .I1(in[84]),
    .O(v1[20])
  );
LUT2  #(
    .INIT(4'h6)
  ) _029_ (
    .I0(in[117]),
    .I1(in[85]),
    .O(v1[21])
  );
LUT2  #(
    .INIT(4'h6)
  ) _030_ (
    .I0(in[118]),
    .I1(in[86]),
    .O(v1[22])
  );
LUT2  #(
    .INIT(4'h6)
  ) _031_ (
    .I0(in[119]),
    .I1(in[87]),
    .O(v1[23])
  );
LUT3  #(
    .INIT(8'h96)
  ) _032_ (
    .I0(in[120]),
    .I1(rcon[0]),
    .I2(in[88]),
    .O(v1[24])
  );
LUT3  #(
    .INIT(8'h96)
  ) _033_ (
    .I0(in[121]),
    .I1(rcon[1]),
    .I2(in[89]),
    .O(v1[25])
  );
LUT3  #(
    .INIT(8'h96)
  ) _034_ (
    .I0(in[122]),
    .I1(rcon[2]),
    .I2(in[90]),
    .O(v1[26])
  );
LUT3  #(
    .INIT(8'h96)
  ) _035_ (
    .I0(in[123]),
    .I1(rcon[3]),
    .I2(in[91]),
    .O(v1[27])
  );
LUT3  #(
    .INIT(8'h96)
  ) _036_ (
    .I0(in[124]),
    .I1(rcon[4]),
    .I2(in[92]),
    .O(v1[28])
  );
LUT3  #(
    .INIT(8'h96)
  ) _037_ (
    .I0(in[125]),
    .I1(rcon[5]),
    .I2(in[93]),
    .O(v1[29])
  );
LUT3  #(
    .INIT(8'h96)
  ) _038_ (
    .I0(in[126]),
    .I1(rcon[6]),
    .I2(in[94]),
    .O(v1[30])
  );
LUT3  #(
    .INIT(8'h96)
  ) _039_ (
    .I0(in[127]),
    .I1(rcon[7]),
    .I2(in[95]),
    .O(v1[31])
  );
LUT3  #(
    .INIT(8'h96)
  ) _040_ (
    .I0(in[96]),
    .I1(in[64]),
    .I2(in[32]),
    .O(v2[0])
  );
LUT3  #(
    .INIT(8'h96)
  ) _041_ (
    .I0(in[97]),
    .I1(in[65]),
    .I2(in[33]),
    .O(v2[1])
  );
LUT3  #(
    .INIT(8'h96)
  ) _042_ (
    .I0(in[98]),
    .I1(in[66]),
    .I2(in[34]),
    .O(v2[2])
  );
LUT3  #(
    .INIT(8'h96)
  ) _043_ (
    .I0(in[99]),
    .I1(in[67]),
    .I2(in[35]),
    .O(v2[3])
  );
LUT3  #(
    .INIT(8'h96)
  ) _044_ (
    .I0(in[100]),
    .I1(in[68]),
    .I2(in[36]),
    .O(v2[4])
  );
LUT3  #(
    .INIT(8'h96)
  ) _045_ (
    .I0(in[101]),
    .I1(in[69]),
    .I2(in[37]),
    .O(v2[5])
  );
LUT3  #(
    .INIT(8'h96)
  ) _046_ (
    .I0(in[102]),
    .I1(in[70]),
    .I2(in[38]),
    .O(v2[6])
  );
LUT3  #(
    .INIT(8'h96)
  ) _047_ (
    .I0(in[103]),
    .I1(in[71]),
    .I2(in[39]),
    .O(v2[7])
  );
LUT3  #(
    .INIT(8'h96)
  ) _048_ (
    .I0(in[104]),
    .I1(in[72]),
    .I2(in[40]),
    .O(v2[8])
  );
LUT3  #(
    .INIT(8'h96)
  ) _049_ (
    .I0(in[105]),
    .I1(in[73]),
    .I2(in[41]),
    .O(v2[9])
  );
LUT3  #(
    .INIT(8'h96)
  ) _050_ (
    .I0(in[106]),
    .I1(in[74]),
    .I2(in[42]),
    .O(v2[10])
  );
LUT3  #(
    .INIT(8'h96)
  ) _051_ (
    .I0(in[107]),
    .I1(in[75]),
    .I2(in[43]),
    .O(v2[11])
  );
LUT3  #(
    .INIT(8'h96)
  ) _052_ (
    .I0(in[108]),
    .I1(in[76]),
    .I2(in[44]),
    .O(v2[12])
  );
LUT3  #(
    .INIT(8'h96)
  ) _053_ (
    .I0(in[109]),
    .I1(in[77]),
    .I2(in[45]),
    .O(v2[13])
  );
LUT3  #(
    .INIT(8'h96)
  ) _054_ (
    .I0(in[110]),
    .I1(in[78]),
    .I2(in[46]),
    .O(v2[14])
  );
LUT3  #(
    .INIT(8'h96)
  ) _055_ (
    .I0(in[111]),
    .I1(in[79]),
    .I2(in[47]),
    .O(v2[15])
  );
LUT3  #(
    .INIT(8'h96)
  ) _056_ (
    .I0(in[112]),
    .I1(in[80]),
    .I2(in[48]),
    .O(v2[16])
  );
LUT3  #(
    .INIT(8'h96)
  ) _057_ (
    .I0(in[113]),
    .I1(in[81]),
    .I2(in[49]),
    .O(v2[17])
  );
LUT3  #(
    .INIT(8'h96)
  ) _058_ (
    .I0(in[114]),
    .I1(in[82]),
    .I2(in[50]),
    .O(v2[18])
  );
LUT3  #(
    .INIT(8'h96)
  ) _059_ (
    .I0(in[115]),
    .I1(in[83]),
    .I2(in[51]),
    .O(v2[19])
  );
LUT3  #(
    .INIT(8'h96)
  ) _060_ (
    .I0(in[116]),
    .I1(in[84]),
    .I2(in[52]),
    .O(v2[20])
  );
LUT3  #(
    .INIT(8'h96)
  ) _061_ (
    .I0(in[117]),
    .I1(in[85]),
    .I2(in[53]),
    .O(v2[21])
  );
LUT3  #(
    .INIT(8'h96)
  ) _062_ (
    .I0(in[118]),
    .I1(in[86]),
    .I2(in[54]),
    .O(v2[22])
  );
LUT3  #(
    .INIT(8'h96)
  ) _063_ (
    .I0(in[119]),
    .I1(in[87]),
    .I2(in[55]),
    .O(v2[23])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _064_ (
    .I0(in[120]),
    .I1(rcon[0]),
    .I2(in[88]),
    .I3(in[56]),
    .O(v2[24])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _065_ (
    .I0(in[121]),
    .I1(rcon[1]),
    .I2(in[89]),
    .I3(in[57]),
    .O(v2[25])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _066_ (
    .I0(in[122]),
    .I1(rcon[2]),
    .I2(in[90]),
    .I3(in[58]),
    .O(v2[26])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _067_ (
    .I0(in[123]),
    .I1(rcon[3]),
    .I2(in[91]),
    .I3(in[59]),
    .O(v2[27])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _068_ (
    .I0(in[124]),
    .I1(rcon[4]),
    .I2(in[92]),
    .I3(in[60]),
    .O(v2[28])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _069_ (
    .I0(in[125]),
    .I1(rcon[5]),
    .I2(in[93]),
    .I3(in[61]),
    .O(v2[29])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _070_ (
    .I0(in[126]),
    .I1(rcon[6]),
    .I2(in[94]),
    .I3(in[62]),
    .O(v2[30])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _071_ (
    .I0(in[127]),
    .I1(rcon[7]),
    .I2(in[95]),
    .I3(in[63]),
    .O(v2[31])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _072_ (
    .I0(in[96]),
    .I1(in[64]),
    .I2(in[32]),
    .I3(in[0]),
    .O(v3[0])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _073_ (
    .I0(in[97]),
    .I1(in[65]),
    .I2(in[33]),
    .I3(in[1]),
    .O(v3[1])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _074_ (
    .I0(in[98]),
    .I1(in[66]),
    .I2(in[34]),
    .I3(in[2]),
    .O(v3[2])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _075_ (
    .I0(in[99]),
    .I1(in[67]),
    .I2(in[35]),
    .I3(in[3]),
    .O(v3[3])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _076_ (
    .I0(in[100]),
    .I1(in[68]),
    .I2(in[36]),
    .I3(in[4]),
    .O(v3[4])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _077_ (
    .I0(in[101]),
    .I1(in[69]),
    .I2(in[37]),
    .I3(in[5]),
    .O(v3[5])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _078_ (
    .I0(in[102]),
    .I1(in[70]),
    .I2(in[38]),
    .I3(in[6]),
    .O(v3[6])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _079_ (
    .I0(in[103]),
    .I1(in[71]),
    .I2(in[39]),
    .I3(in[7]),
    .O(v3[7])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _080_ (
    .I0(in[104]),
    .I1(in[72]),
    .I2(in[40]),
    .I3(in[8]),
    .O(v3[8])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _081_ (
    .I0(in[105]),
    .I1(in[73]),
    .I2(in[41]),
    .I3(in[9]),
    .O(v3[9])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _082_ (
    .I0(in[106]),
    .I1(in[74]),
    .I2(in[42]),
    .I3(in[10]),
    .O(v3[10])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _083_ (
    .I0(in[107]),
    .I1(in[75]),
    .I2(in[43]),
    .I3(in[11]),
    .O(v3[11])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _084_ (
    .I0(in[108]),
    .I1(in[76]),
    .I2(in[44]),
    .I3(in[12]),
    .O(v3[12])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _085_ (
    .I0(in[109]),
    .I1(in[77]),
    .I2(in[45]),
    .I3(in[13]),
    .O(v3[13])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _086_ (
    .I0(in[110]),
    .I1(in[78]),
    .I2(in[46]),
    .I3(in[14]),
    .O(v3[14])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _087_ (
    .I0(in[111]),
    .I1(in[79]),
    .I2(in[47]),
    .I3(in[15]),
    .O(v3[15])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _088_ (
    .I0(in[112]),
    .I1(in[80]),
    .I2(in[48]),
    .I3(in[16]),
    .O(v3[16])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _089_ (
    .I0(in[113]),
    .I1(in[81]),
    .I2(in[49]),
    .I3(in[17]),
    .O(v3[17])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _090_ (
    .I0(in[114]),
    .I1(in[82]),
    .I2(in[50]),
    .I3(in[18]),
    .O(v3[18])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _091_ (
    .I0(in[115]),
    .I1(in[83]),
    .I2(in[51]),
    .I3(in[19]),
    .O(v3[19])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _092_ (
    .I0(in[116]),
    .I1(in[84]),
    .I2(in[52]),
    .I3(in[20]),
    .O(v3[20])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _093_ (
    .I0(in[117]),
    .I1(in[85]),
    .I2(in[53]),
    .I3(in[21]),
    .O(v3[21])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _094_ (
    .I0(in[118]),
    .I1(in[86]),
    .I2(in[54]),
    .I3(in[22]),
    .O(v3[22])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _095_ (
    .I0(in[119]),
    .I1(in[87]),
    .I2(in[55]),
    .I3(in[23]),
    .O(v3[23])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _096_ (
    .I0(in[120]),
    .I1(rcon[0]),
    .I2(in[88]),
    .I3(in[56]),
    .I4(in[24]),
    .O(v3[24])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _097_ (
    .I0(in[121]),
    .I1(rcon[1]),
    .I2(in[89]),
    .I3(in[57]),
    .I4(in[25]),
    .O(v3[25])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _098_ (
    .I0(in[122]),
    .I1(rcon[2]),
    .I2(in[90]),
    .I3(in[58]),
    .I4(in[26]),
    .O(v3[26])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _099_ (
    .I0(in[123]),
    .I1(rcon[3]),
    .I2(in[91]),
    .I3(in[59]),
    .I4(in[27]),
    .O(v3[27])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _100_ (
    .I0(in[124]),
    .I1(rcon[4]),
    .I2(in[92]),
    .I3(in[60]),
    .I4(in[28]),
    .O(v3[28])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _101_ (
    .I0(in[125]),
    .I1(rcon[5]),
    .I2(in[93]),
    .I3(in[61]),
    .I4(in[29]),
    .O(v3[29])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _102_ (
    .I0(in[126]),
    .I1(rcon[6]),
    .I2(in[94]),
    .I3(in[62]),
    .I4(in[30]),
    .O(v3[30])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _103_ (
    .I0(in[127]),
    .I1(rcon[7]),
    .I2(in[95]),
    .I3(in[63]),
    .I4(in[31]),
    .O(v3[31])
  );
LUT2  #(
    .INIT(4'h6)
  ) _104_ (
    .I0(k0a[0]),
    .I1(k4a[0]),
    .O(k0b[0])
  );
LUT2  #(
    .INIT(4'h6)
  ) _105_ (
    .I0(k0a[1]),
    .I1(k4a[1]),
    .O(k0b[1])
  );
LUT2  #(
    .INIT(4'h6)
  ) _106_ (
    .I0(k0a[2]),
    .I1(k4a[2]),
    .O(k0b[2])
  );
LUT2  #(
    .INIT(4'h6)
  ) _107_ (
    .I0(k0a[3]),
    .I1(k4a[3]),
    .O(k0b[3])
  );
LUT2  #(
    .INIT(4'h6)
  ) _108_ (
    .I0(k0a[4]),
    .I1(k4a[4]),
    .O(k0b[4])
  );
LUT2  #(
    .INIT(4'h6)
  ) _109_ (
    .I0(k0a[5]),
    .I1(k4a[5]),
    .O(k0b[5])
  );
LUT2  #(
    .INIT(4'h6)
  ) _110_ (
    .I0(k0a[6]),
    .I1(k4a[6]),
    .O(k0b[6])
  );
LUT2  #(
    .INIT(4'h6)
  ) _111_ (
    .I0(k0a[7]),
    .I1(k4a[7]),
    .O(k0b[7])
  );
LUT2  #(
    .INIT(4'h6)
  ) _112_ (
    .I0(k0a[8]),
    .I1(k4a[8]),
    .O(k0b[8])
  );
LUT2  #(
    .INIT(4'h6)
  ) _113_ (
    .I0(k0a[9]),
    .I1(k4a[9]),
    .O(k0b[9])
  );
LUT2  #(
    .INIT(4'h6)
  ) _114_ (
    .I0(k0a[10]),
    .I1(k4a[10]),
    .O(k0b[10])
  );
LUT2  #(
    .INIT(4'h6)
  ) _115_ (
    .I0(k0a[11]),
    .I1(k4a[11]),
    .O(k0b[11])
  );
LUT2  #(
    .INIT(4'h6)
  ) _116_ (
    .I0(k0a[12]),
    .I1(k4a[12]),
    .O(k0b[12])
  );
LUT2  #(
    .INIT(4'h6)
  ) _117_ (
    .I0(k0a[13]),
    .I1(k4a[13]),
    .O(k0b[13])
  );
LUT2  #(
    .INIT(4'h6)
  ) _118_ (
    .I0(k0a[14]),
    .I1(k4a[14]),
    .O(k0b[14])
  );
LUT2  #(
    .INIT(4'h6)
  ) _119_ (
    .I0(k0a[15]),
    .I1(k4a[15]),
    .O(k0b[15])
  );
LUT2  #(
    .INIT(4'h6)
  ) _120_ (
    .I0(k0a[16]),
    .I1(k4a[16]),
    .O(k0b[16])
  );
LUT2  #(
    .INIT(4'h6)
  ) _121_ (
    .I0(k0a[17]),
    .I1(k4a[17]),
    .O(k0b[17])
  );
LUT2  #(
    .INIT(4'h6)
  ) _122_ (
    .I0(k0a[18]),
    .I1(k4a[18]),
    .O(k0b[18])
  );
LUT2  #(
    .INIT(4'h6)
  ) _123_ (
    .I0(k0a[19]),
    .I1(k4a[19]),
    .O(k0b[19])
  );
LUT2  #(
    .INIT(4'h6)
  ) _124_ (
    .I0(k0a[20]),
    .I1(k4a[20]),
    .O(k0b[20])
  );
LUT2  #(
    .INIT(4'h6)
  ) _125_ (
    .I0(k0a[21]),
    .I1(k4a[21]),
    .O(k0b[21])
  );
LUT2  #(
    .INIT(4'h6)
  ) _126_ (
    .I0(k0a[22]),
    .I1(k4a[22]),
    .O(k0b[22])
  );
LUT2  #(
    .INIT(4'h6)
  ) _127_ (
    .I0(k0a[23]),
    .I1(k4a[23]),
    .O(k0b[23])
  );
LUT2  #(
    .INIT(4'h6)
  ) _128_ (
    .I0(k0a[24]),
    .I1(k4a[24]),
    .O(k0b[24])
  );
LUT2  #(
    .INIT(4'h6)
  ) _129_ (
    .I0(k0a[25]),
    .I1(k4a[25]),
    .O(k0b[25])
  );
LUT2  #(
    .INIT(4'h6)
  ) _130_ (
    .I0(k0a[26]),
    .I1(k4a[26]),
    .O(k0b[26])
  );
LUT2  #(
    .INIT(4'h6)
  ) _131_ (
    .I0(k0a[27]),
    .I1(k4a[27]),
    .O(k0b[27])
  );
LUT2  #(
    .INIT(4'h6)
  ) _132_ (
    .I0(k0a[28]),
    .I1(k4a[28]),
    .O(k0b[28])
  );
LUT2  #(
    .INIT(4'h6)
  ) _133_ (
    .I0(k0a[29]),
    .I1(k4a[29]),
    .O(k0b[29])
  );
LUT2  #(
    .INIT(4'h6)
  ) _134_ (
    .I0(k0a[30]),
    .I1(k4a[30]),
    .O(k0b[30])
  );
LUT2  #(
    .INIT(4'h6)
  ) _135_ (
    .I0(k0a[31]),
    .I1(k4a[31]),
    .O(k0b[31])
  );
LUT2  #(
    .INIT(4'h6)
  ) _136_ (
    .I0(k4a[0]),
    .I1(k1a[0]),
    .O(k1b[0])
  );
LUT2  #(
    .INIT(4'h6)
  ) _137_ (
    .I0(k4a[1]),
    .I1(k1a[1]),
    .O(k1b[1])
  );
LUT2  #(
    .INIT(4'h6)
  ) _138_ (
    .I0(k4a[2]),
    .I1(k1a[2]),
    .O(k1b[2])
  );
LUT2  #(
    .INIT(4'h6)
  ) _139_ (
    .I0(k4a[3]),
    .I1(k1a[3]),
    .O(k1b[3])
  );
LUT2  #(
    .INIT(4'h6)
  ) _140_ (
    .I0(k4a[4]),
    .I1(k1a[4]),
    .O(k1b[4])
  );
LUT2  #(
    .INIT(4'h6)
  ) _141_ (
    .I0(k4a[5]),
    .I1(k1a[5]),
    .O(k1b[5])
  );
LUT2  #(
    .INIT(4'h6)
  ) _142_ (
    .I0(k4a[6]),
    .I1(k1a[6]),
    .O(k1b[6])
  );
LUT2  #(
    .INIT(4'h6)
  ) _143_ (
    .I0(k4a[7]),
    .I1(k1a[7]),
    .O(k1b[7])
  );
LUT2  #(
    .INIT(4'h6)
  ) _144_ (
    .I0(k4a[8]),
    .I1(k1a[8]),
    .O(k1b[8])
  );
LUT2  #(
    .INIT(4'h6)
  ) _145_ (
    .I0(k4a[9]),
    .I1(k1a[9]),
    .O(k1b[9])
  );
LUT2  #(
    .INIT(4'h6)
  ) _146_ (
    .I0(k4a[10]),
    .I1(k1a[10]),
    .O(k1b[10])
  );
LUT2  #(
    .INIT(4'h6)
  ) _147_ (
    .I0(k4a[11]),
    .I1(k1a[11]),
    .O(k1b[11])
  );
LUT2  #(
    .INIT(4'h6)
  ) _148_ (
    .I0(k4a[12]),
    .I1(k1a[12]),
    .O(k1b[12])
  );
LUT2  #(
    .INIT(4'h6)
  ) _149_ (
    .I0(k4a[13]),
    .I1(k1a[13]),
    .O(k1b[13])
  );
LUT2  #(
    .INIT(4'h6)
  ) _150_ (
    .I0(k4a[14]),
    .I1(k1a[14]),
    .O(k1b[14])
  );
LUT2  #(
    .INIT(4'h6)
  ) _151_ (
    .I0(k4a[15]),
    .I1(k1a[15]),
    .O(k1b[15])
  );
LUT2  #(
    .INIT(4'h6)
  ) _152_ (
    .I0(k4a[16]),
    .I1(k1a[16]),
    .O(k1b[16])
  );
LUT2  #(
    .INIT(4'h6)
  ) _153_ (
    .I0(k4a[17]),
    .I1(k1a[17]),
    .O(k1b[17])
  );
LUT2  #(
    .INIT(4'h6)
  ) _154_ (
    .I0(k4a[18]),
    .I1(k1a[18]),
    .O(k1b[18])
  );
LUT2  #(
    .INIT(4'h6)
  ) _155_ (
    .I0(k4a[19]),
    .I1(k1a[19]),
    .O(k1b[19])
  );
LUT2  #(
    .INIT(4'h6)
  ) _156_ (
    .I0(k4a[20]),
    .I1(k1a[20]),
    .O(k1b[20])
  );
LUT2  #(
    .INIT(4'h6)
  ) _157_ (
    .I0(k4a[21]),
    .I1(k1a[21]),
    .O(k1b[21])
  );
LUT2  #(
    .INIT(4'h6)
  ) _158_ (
    .I0(k4a[22]),
    .I1(k1a[22]),
    .O(k1b[22])
  );
LUT2  #(
    .INIT(4'h6)
  ) _159_ (
    .I0(k4a[23]),
    .I1(k1a[23]),
    .O(k1b[23])
  );
LUT2  #(
    .INIT(4'h6)
  ) _160_ (
    .I0(k4a[24]),
    .I1(k1a[24]),
    .O(k1b[24])
  );
LUT2  #(
    .INIT(4'h6)
  ) _161_ (
    .I0(k4a[25]),
    .I1(k1a[25]),
    .O(k1b[25])
  );
LUT2  #(
    .INIT(4'h6)
  ) _162_ (
    .I0(k4a[26]),
    .I1(k1a[26]),
    .O(k1b[26])
  );
LUT2  #(
    .INIT(4'h6)
  ) _163_ (
    .I0(k4a[27]),
    .I1(k1a[27]),
    .O(k1b[27])
  );
LUT2  #(
    .INIT(4'h6)
  ) _164_ (
    .I0(k4a[28]),
    .I1(k1a[28]),
    .O(k1b[28])
  );
LUT2  #(
    .INIT(4'h6)
  ) _165_ (
    .I0(k4a[29]),
    .I1(k1a[29]),
    .O(k1b[29])
  );
LUT2  #(
    .INIT(4'h6)
  ) _166_ (
    .I0(k4a[30]),
    .I1(k1a[30]),
    .O(k1b[30])
  );
LUT2  #(
    .INIT(4'h6)
  ) _167_ (
    .I0(k4a[31]),
    .I1(k1a[31]),
    .O(k1b[31])
  );
LUT2  #(
    .INIT(4'h6)
  ) _168_ (
    .I0(k4a[0]),
    .I1(k2a[0]),
    .O(k2b[0])
  );
LUT2  #(
    .INIT(4'h6)
  ) _169_ (
    .I0(k4a[1]),
    .I1(k2a[1]),
    .O(k2b[1])
  );
LUT2  #(
    .INIT(4'h6)
  ) _170_ (
    .I0(k4a[2]),
    .I1(k2a[2]),
    .O(k2b[2])
  );
LUT2  #(
    .INIT(4'h6)
  ) _171_ (
    .I0(k4a[3]),
    .I1(k2a[3]),
    .O(k2b[3])
  );
LUT2  #(
    .INIT(4'h6)
  ) _172_ (
    .I0(k4a[4]),
    .I1(k2a[4]),
    .O(k2b[4])
  );
LUT2  #(
    .INIT(4'h6)
  ) _173_ (
    .I0(k4a[5]),
    .I1(k2a[5]),
    .O(k2b[5])
  );
LUT2  #(
    .INIT(4'h6)
  ) _174_ (
    .I0(k4a[6]),
    .I1(k2a[6]),
    .O(k2b[6])
  );
LUT2  #(
    .INIT(4'h6)
  ) _175_ (
    .I0(k4a[7]),
    .I1(k2a[7]),
    .O(k2b[7])
  );
LUT2  #(
    .INIT(4'h6)
  ) _176_ (
    .I0(k4a[8]),
    .I1(k2a[8]),
    .O(k2b[8])
  );
LUT2  #(
    .INIT(4'h6)
  ) _177_ (
    .I0(k4a[9]),
    .I1(k2a[9]),
    .O(k2b[9])
  );
LUT2  #(
    .INIT(4'h6)
  ) _178_ (
    .I0(k4a[10]),
    .I1(k2a[10]),
    .O(k2b[10])
  );
LUT2  #(
    .INIT(4'h6)
  ) _179_ (
    .I0(k4a[11]),
    .I1(k2a[11]),
    .O(k2b[11])
  );
LUT2  #(
    .INIT(4'h6)
  ) _180_ (
    .I0(k4a[12]),
    .I1(k2a[12]),
    .O(k2b[12])
  );
LUT2  #(
    .INIT(4'h6)
  ) _181_ (
    .I0(k4a[13]),
    .I1(k2a[13]),
    .O(k2b[13])
  );
LUT2  #(
    .INIT(4'h6)
  ) _182_ (
    .I0(k4a[14]),
    .I1(k2a[14]),
    .O(k2b[14])
  );
LUT2  #(
    .INIT(4'h6)
  ) _183_ (
    .I0(k4a[15]),
    .I1(k2a[15]),
    .O(k2b[15])
  );
LUT2  #(
    .INIT(4'h6)
  ) _184_ (
    .I0(k4a[16]),
    .I1(k2a[16]),
    .O(k2b[16])
  );
LUT2  #(
    .INIT(4'h6)
  ) _185_ (
    .I0(k4a[17]),
    .I1(k2a[17]),
    .O(k2b[17])
  );
LUT2  #(
    .INIT(4'h6)
  ) _186_ (
    .I0(k4a[18]),
    .I1(k2a[18]),
    .O(k2b[18])
  );
LUT2  #(
    .INIT(4'h6)
  ) _187_ (
    .I0(k4a[19]),
    .I1(k2a[19]),
    .O(k2b[19])
  );
LUT2  #(
    .INIT(4'h6)
  ) _188_ (
    .I0(k4a[20]),
    .I1(k2a[20]),
    .O(k2b[20])
  );
LUT2  #(
    .INIT(4'h6)
  ) _189_ (
    .I0(k4a[21]),
    .I1(k2a[21]),
    .O(k2b[21])
  );
LUT2  #(
    .INIT(4'h6)
  ) _190_ (
    .I0(k4a[22]),
    .I1(k2a[22]),
    .O(k2b[22])
  );
LUT2  #(
    .INIT(4'h6)
  ) _191_ (
    .I0(k4a[23]),
    .I1(k2a[23]),
    .O(k2b[23])
  );
LUT2  #(
    .INIT(4'h6)
  ) _192_ (
    .I0(k4a[24]),
    .I1(k2a[24]),
    .O(k2b[24])
  );
LUT2  #(
    .INIT(4'h6)
  ) _193_ (
    .I0(k4a[25]),
    .I1(k2a[25]),
    .O(k2b[25])
  );
LUT2  #(
    .INIT(4'h6)
  ) _194_ (
    .I0(k4a[26]),
    .I1(k2a[26]),
    .O(k2b[26])
  );
LUT2  #(
    .INIT(4'h6)
  ) _195_ (
    .I0(k4a[27]),
    .I1(k2a[27]),
    .O(k2b[27])
  );
LUT2  #(
    .INIT(4'h6)
  ) _196_ (
    .I0(k4a[28]),
    .I1(k2a[28]),
    .O(k2b[28])
  );
LUT2  #(
    .INIT(4'h6)
  ) _197_ (
    .I0(k4a[29]),
    .I1(k2a[29]),
    .O(k2b[29])
  );
LUT2  #(
    .INIT(4'h6)
  ) _198_ (
    .I0(k4a[30]),
    .I1(k2a[30]),
    .O(k2b[30])
  );
LUT2  #(
    .INIT(4'h6)
  ) _199_ (
    .I0(k4a[31]),
    .I1(k2a[31]),
    .O(k2b[31])
  );
LUT2  #(
    .INIT(4'h6)
  ) _200_ (
    .I0(k4a[0]),
    .I1(k3a[0]),
    .O(k3b[0])
  );
LUT2  #(
    .INIT(4'h6)
  ) _201_ (
    .I0(k4a[1]),
    .I1(k3a[1]),
    .O(k3b[1])
  );
LUT2  #(
    .INIT(4'h6)
  ) _202_ (
    .I0(k4a[2]),
    .I1(k3a[2]),
    .O(k3b[2])
  );
LUT2  #(
    .INIT(4'h6)
  ) _203_ (
    .I0(k4a[3]),
    .I1(k3a[3]),
    .O(k3b[3])
  );
LUT2  #(
    .INIT(4'h6)
  ) _204_ (
    .I0(k4a[4]),
    .I1(k3a[4]),
    .O(k3b[4])
  );
LUT2  #(
    .INIT(4'h6)
  ) _205_ (
    .I0(k4a[5]),
    .I1(k3a[5]),
    .O(k3b[5])
  );
LUT2  #(
    .INIT(4'h6)
  ) _206_ (
    .I0(k4a[6]),
    .I1(k3a[6]),
    .O(k3b[6])
  );
LUT2  #(
    .INIT(4'h6)
  ) _207_ (
    .I0(k4a[7]),
    .I1(k3a[7]),
    .O(k3b[7])
  );
LUT2  #(
    .INIT(4'h6)
  ) _208_ (
    .I0(k4a[8]),
    .I1(k3a[8]),
    .O(k3b[8])
  );
LUT2  #(
    .INIT(4'h6)
  ) _209_ (
    .I0(k4a[9]),
    .I1(k3a[9]),
    .O(k3b[9])
  );
LUT2  #(
    .INIT(4'h6)
  ) _210_ (
    .I0(k4a[10]),
    .I1(k3a[10]),
    .O(k3b[10])
  );
LUT2  #(
    .INIT(4'h6)
  ) _211_ (
    .I0(k4a[11]),
    .I1(k3a[11]),
    .O(k3b[11])
  );
LUT2  #(
    .INIT(4'h6)
  ) _212_ (
    .I0(k4a[12]),
    .I1(k3a[12]),
    .O(k3b[12])
  );
LUT2  #(
    .INIT(4'h6)
  ) _213_ (
    .I0(k4a[13]),
    .I1(k3a[13]),
    .O(k3b[13])
  );
LUT2  #(
    .INIT(4'h6)
  ) _214_ (
    .I0(k4a[14]),
    .I1(k3a[14]),
    .O(k3b[14])
  );
LUT2  #(
    .INIT(4'h6)
  ) _215_ (
    .I0(k4a[15]),
    .I1(k3a[15]),
    .O(k3b[15])
  );
LUT2  #(
    .INIT(4'h6)
  ) _216_ (
    .I0(k4a[16]),
    .I1(k3a[16]),
    .O(k3b[16])
  );
LUT2  #(
    .INIT(4'h6)
  ) _217_ (
    .I0(k4a[17]),
    .I1(k3a[17]),
    .O(k3b[17])
  );
LUT2  #(
    .INIT(4'h6)
  ) _218_ (
    .I0(k4a[18]),
    .I1(k3a[18]),
    .O(k3b[18])
  );
LUT2  #(
    .INIT(4'h6)
  ) _219_ (
    .I0(k4a[19]),
    .I1(k3a[19]),
    .O(k3b[19])
  );
LUT2  #(
    .INIT(4'h6)
  ) _220_ (
    .I0(k4a[20]),
    .I1(k3a[20]),
    .O(k3b[20])
  );
LUT2  #(
    .INIT(4'h6)
  ) _221_ (
    .I0(k4a[21]),
    .I1(k3a[21]),
    .O(k3b[21])
  );
LUT2  #(
    .INIT(4'h6)
  ) _222_ (
    .I0(k4a[22]),
    .I1(k3a[22]),
    .O(k3b[22])
  );
LUT2  #(
    .INIT(4'h6)
  ) _223_ (
    .I0(k4a[23]),
    .I1(k3a[23]),
    .O(k3b[23])
  );
LUT2  #(
    .INIT(4'h6)
  ) _224_ (
    .I0(k4a[24]),
    .I1(k3a[24]),
    .O(k3b[24])
  );
LUT2  #(
    .INIT(4'h6)
  ) _225_ (
    .I0(k4a[25]),
    .I1(k3a[25]),
    .O(k3b[25])
  );
LUT2  #(
    .INIT(4'h6)
  ) _226_ (
    .I0(k4a[26]),
    .I1(k3a[26]),
    .O(k3b[26])
  );
LUT2  #(
    .INIT(4'h6)
  ) _227_ (
    .I0(k4a[27]),
    .I1(k3a[27]),
    .O(k3b[27])
  );
LUT2  #(
    .INIT(4'h6)
  ) _228_ (
    .I0(k4a[28]),
    .I1(k3a[28]),
    .O(k3b[28])
  );
LUT2  #(
    .INIT(4'h6)
  ) _229_ (
    .I0(k4a[29]),
    .I1(k3a[29]),
    .O(k3b[29])
  );
LUT2  #(
    .INIT(4'h6)
  ) _230_ (
    .I0(k4a[30]),
    .I1(k3a[30]),
    .O(k3b[30])
  );
LUT2  #(
    .INIT(4'h6)
  ) _231_ (
    .I0(k4a[31]),
    .I1(k3a[31]),
    .O(k3b[31])
  );
FDRE  #(
    .INIT(1'hx)
  ) _232_ (
    .C(clk),
    .CE(1'h1),
    .D(k3b[0]),
    .Q(out_1[0]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _233_ (
    .C(clk),
    .CE(1'h1),
    .D(k3b[1]),
    .Q(out_1[1]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _234_ (
    .C(clk),
    .CE(1'h1),
    .D(k3b[2]),
    .Q(out_1[2]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _235_ (
    .C(clk),
    .CE(1'h1),
    .D(k3b[3]),
    .Q(out_1[3]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _236_ (
    .C(clk),
    .CE(1'h1),
    .D(k3b[4]),
    .Q(out_1[4]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _237_ (
    .C(clk),
    .CE(1'h1),
    .D(k3b[5]),
    .Q(out_1[5]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _238_ (
    .C(clk),
    .CE(1'h1),
    .D(k3b[6]),
    .Q(out_1[6]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _239_ (
    .C(clk),
    .CE(1'h1),
    .D(k3b[7]),
    .Q(out_1[7]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _240_ (
    .C(clk),
    .CE(1'h1),
    .D(k3b[8]),
    .Q(out_1[8]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _241_ (
    .C(clk),
    .CE(1'h1),
    .D(k3b[9]),
    .Q(out_1[9]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _242_ (
    .C(clk),
    .CE(1'h1),
    .D(k3b[10]),
    .Q(out_1[10]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _243_ (
    .C(clk),
    .CE(1'h1),
    .D(k3b[11]),
    .Q(out_1[11]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _244_ (
    .C(clk),
    .CE(1'h1),
    .D(k3b[12]),
    .Q(out_1[12]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _245_ (
    .C(clk),
    .CE(1'h1),
    .D(k3b[13]),
    .Q(out_1[13]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _246_ (
    .C(clk),
    .CE(1'h1),
    .D(k3b[14]),
    .Q(out_1[14]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _247_ (
    .C(clk),
    .CE(1'h1),
    .D(k3b[15]),
    .Q(out_1[15]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _248_ (
    .C(clk),
    .CE(1'h1),
    .D(k3b[16]),
    .Q(out_1[16]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _249_ (
    .C(clk),
    .CE(1'h1),
    .D(k3b[17]),
    .Q(out_1[17]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _250_ (
    .C(clk),
    .CE(1'h1),
    .D(k3b[18]),
    .Q(out_1[18]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _251_ (
    .C(clk),
    .CE(1'h1),
    .D(k3b[19]),
    .Q(out_1[19]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _252_ (
    .C(clk),
    .CE(1'h1),
    .D(k3b[20]),
    .Q(out_1[20]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _253_ (
    .C(clk),
    .CE(1'h1),
    .D(k3b[21]),
    .Q(out_1[21]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _254_ (
    .C(clk),
    .CE(1'h1),
    .D(k3b[22]),
    .Q(out_1[22]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _255_ (
    .C(clk),
    .CE(1'h1),
    .D(k3b[23]),
    .Q(out_1[23]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _256_ (
    .C(clk),
    .CE(1'h1),
    .D(k3b[24]),
    .Q(out_1[24]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _257_ (
    .C(clk),
    .CE(1'h1),
    .D(k3b[25]),
    .Q(out_1[25]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _258_ (
    .C(clk),
    .CE(1'h1),
    .D(k3b[26]),
    .Q(out_1[26]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _259_ (
    .C(clk),
    .CE(1'h1),
    .D(k3b[27]),
    .Q(out_1[27]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _260_ (
    .C(clk),
    .CE(1'h1),
    .D(k3b[28]),
    .Q(out_1[28]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _261_ (
    .C(clk),
    .CE(1'h1),
    .D(k3b[29]),
    .Q(out_1[29]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _262_ (
    .C(clk),
    .CE(1'h1),
    .D(k3b[30]),
    .Q(out_1[30]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _263_ (
    .C(clk),
    .CE(1'h1),
    .D(k3b[31]),
    .Q(out_1[31]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _264_ (
    .C(clk),
    .CE(1'h1),
    .D(k2b[0]),
    .Q(out_1[32]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _265_ (
    .C(clk),
    .CE(1'h1),
    .D(k2b[1]),
    .Q(out_1[33]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _266_ (
    .C(clk),
    .CE(1'h1),
    .D(k2b[2]),
    .Q(out_1[34]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _267_ (
    .C(clk),
    .CE(1'h1),
    .D(k2b[3]),
    .Q(out_1[35]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _268_ (
    .C(clk),
    .CE(1'h1),
    .D(k2b[4]),
    .Q(out_1[36]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _269_ (
    .C(clk),
    .CE(1'h1),
    .D(k2b[5]),
    .Q(out_1[37]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _270_ (
    .C(clk),
    .CE(1'h1),
    .D(k2b[6]),
    .Q(out_1[38]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _271_ (
    .C(clk),
    .CE(1'h1),
    .D(k2b[7]),
    .Q(out_1[39]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _272_ (
    .C(clk),
    .CE(1'h1),
    .D(k2b[8]),
    .Q(out_1[40]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _273_ (
    .C(clk),
    .CE(1'h1),
    .D(k2b[9]),
    .Q(out_1[41]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _274_ (
    .C(clk),
    .CE(1'h1),
    .D(k2b[10]),
    .Q(out_1[42]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _275_ (
    .C(clk),
    .CE(1'h1),
    .D(k2b[11]),
    .Q(out_1[43]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _276_ (
    .C(clk),
    .CE(1'h1),
    .D(k2b[12]),
    .Q(out_1[44]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _277_ (
    .C(clk),
    .CE(1'h1),
    .D(k2b[13]),
    .Q(out_1[45]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _278_ (
    .C(clk),
    .CE(1'h1),
    .D(k2b[14]),
    .Q(out_1[46]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _279_ (
    .C(clk),
    .CE(1'h1),
    .D(k2b[15]),
    .Q(out_1[47]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _280_ (
    .C(clk),
    .CE(1'h1),
    .D(k2b[16]),
    .Q(out_1[48]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _281_ (
    .C(clk),
    .CE(1'h1),
    .D(k2b[17]),
    .Q(out_1[49]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _282_ (
    .C(clk),
    .CE(1'h1),
    .D(k2b[18]),
    .Q(out_1[50]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _283_ (
    .C(clk),
    .CE(1'h1),
    .D(k2b[19]),
    .Q(out_1[51]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _284_ (
    .C(clk),
    .CE(1'h1),
    .D(k2b[20]),
    .Q(out_1[52]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _285_ (
    .C(clk),
    .CE(1'h1),
    .D(k2b[21]),
    .Q(out_1[53]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _286_ (
    .C(clk),
    .CE(1'h1),
    .D(k2b[22]),
    .Q(out_1[54]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _287_ (
    .C(clk),
    .CE(1'h1),
    .D(k2b[23]),
    .Q(out_1[55]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _288_ (
    .C(clk),
    .CE(1'h1),
    .D(k2b[24]),
    .Q(out_1[56]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _289_ (
    .C(clk),
    .CE(1'h1),
    .D(k2b[25]),
    .Q(out_1[57]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _290_ (
    .C(clk),
    .CE(1'h1),
    .D(k2b[26]),
    .Q(out_1[58]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _291_ (
    .C(clk),
    .CE(1'h1),
    .D(k2b[27]),
    .Q(out_1[59]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _292_ (
    .C(clk),
    .CE(1'h1),
    .D(k2b[28]),
    .Q(out_1[60]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _293_ (
    .C(clk),
    .CE(1'h1),
    .D(k2b[29]),
    .Q(out_1[61]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _294_ (
    .C(clk),
    .CE(1'h1),
    .D(k2b[30]),
    .Q(out_1[62]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _295_ (
    .C(clk),
    .CE(1'h1),
    .D(k2b[31]),
    .Q(out_1[63]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _296_ (
    .C(clk),
    .CE(1'h1),
    .D(k1b[0]),
    .Q(out_1[64]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _297_ (
    .C(clk),
    .CE(1'h1),
    .D(k1b[1]),
    .Q(out_1[65]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _298_ (
    .C(clk),
    .CE(1'h1),
    .D(k1b[2]),
    .Q(out_1[66]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _299_ (
    .C(clk),
    .CE(1'h1),
    .D(k1b[3]),
    .Q(out_1[67]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _300_ (
    .C(clk),
    .CE(1'h1),
    .D(k1b[4]),
    .Q(out_1[68]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _301_ (
    .C(clk),
    .CE(1'h1),
    .D(k1b[5]),
    .Q(out_1[69]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _302_ (
    .C(clk),
    .CE(1'h1),
    .D(k1b[6]),
    .Q(out_1[70]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _303_ (
    .C(clk),
    .CE(1'h1),
    .D(k1b[7]),
    .Q(out_1[71]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _304_ (
    .C(clk),
    .CE(1'h1),
    .D(k1b[8]),
    .Q(out_1[72]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _305_ (
    .C(clk),
    .CE(1'h1),
    .D(k1b[9]),
    .Q(out_1[73]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _306_ (
    .C(clk),
    .CE(1'h1),
    .D(k1b[10]),
    .Q(out_1[74]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _307_ (
    .C(clk),
    .CE(1'h1),
    .D(k1b[11]),
    .Q(out_1[75]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _308_ (
    .C(clk),
    .CE(1'h1),
    .D(k1b[12]),
    .Q(out_1[76]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _309_ (
    .C(clk),
    .CE(1'h1),
    .D(k1b[13]),
    .Q(out_1[77]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _310_ (
    .C(clk),
    .CE(1'h1),
    .D(k1b[14]),
    .Q(out_1[78]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _311_ (
    .C(clk),
    .CE(1'h1),
    .D(k1b[15]),
    .Q(out_1[79]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _312_ (
    .C(clk),
    .CE(1'h1),
    .D(k1b[16]),
    .Q(out_1[80]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _313_ (
    .C(clk),
    .CE(1'h1),
    .D(k1b[17]),
    .Q(out_1[81]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _314_ (
    .C(clk),
    .CE(1'h1),
    .D(k1b[18]),
    .Q(out_1[82]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _315_ (
    .C(clk),
    .CE(1'h1),
    .D(k1b[19]),
    .Q(out_1[83]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _316_ (
    .C(clk),
    .CE(1'h1),
    .D(k1b[20]),
    .Q(out_1[84]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _317_ (
    .C(clk),
    .CE(1'h1),
    .D(k1b[21]),
    .Q(out_1[85]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _318_ (
    .C(clk),
    .CE(1'h1),
    .D(k1b[22]),
    .Q(out_1[86]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _319_ (
    .C(clk),
    .CE(1'h1),
    .D(k1b[23]),
    .Q(out_1[87]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _320_ (
    .C(clk),
    .CE(1'h1),
    .D(k1b[24]),
    .Q(out_1[88]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _321_ (
    .C(clk),
    .CE(1'h1),
    .D(k1b[25]),
    .Q(out_1[89]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _322_ (
    .C(clk),
    .CE(1'h1),
    .D(k1b[26]),
    .Q(out_1[90]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _323_ (
    .C(clk),
    .CE(1'h1),
    .D(k1b[27]),
    .Q(out_1[91]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _324_ (
    .C(clk),
    .CE(1'h1),
    .D(k1b[28]),
    .Q(out_1[92]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _325_ (
    .C(clk),
    .CE(1'h1),
    .D(k1b[29]),
    .Q(out_1[93]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _326_ (
    .C(clk),
    .CE(1'h1),
    .D(k1b[30]),
    .Q(out_1[94]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _327_ (
    .C(clk),
    .CE(1'h1),
    .D(k1b[31]),
    .Q(out_1[95]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _328_ (
    .C(clk),
    .CE(1'h1),
    .D(k0b[0]),
    .Q(out_1[96]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _329_ (
    .C(clk),
    .CE(1'h1),
    .D(k0b[1]),
    .Q(out_1[97]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _330_ (
    .C(clk),
    .CE(1'h1),
    .D(k0b[2]),
    .Q(out_1[98]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _331_ (
    .C(clk),
    .CE(1'h1),
    .D(k0b[3]),
    .Q(out_1[99]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _332_ (
    .C(clk),
    .CE(1'h1),
    .D(k0b[4]),
    .Q(out_1[100]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _333_ (
    .C(clk),
    .CE(1'h1),
    .D(k0b[5]),
    .Q(out_1[101]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _334_ (
    .C(clk),
    .CE(1'h1),
    .D(k0b[6]),
    .Q(out_1[102]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _335_ (
    .C(clk),
    .CE(1'h1),
    .D(k0b[7]),
    .Q(out_1[103]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _336_ (
    .C(clk),
    .CE(1'h1),
    .D(k0b[8]),
    .Q(out_1[104]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _337_ (
    .C(clk),
    .CE(1'h1),
    .D(k0b[9]),
    .Q(out_1[105]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _338_ (
    .C(clk),
    .CE(1'h1),
    .D(k0b[10]),
    .Q(out_1[106]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _339_ (
    .C(clk),
    .CE(1'h1),
    .D(k0b[11]),
    .Q(out_1[107]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _340_ (
    .C(clk),
    .CE(1'h1),
    .D(k0b[12]),
    .Q(out_1[108]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _341_ (
    .C(clk),
    .CE(1'h1),
    .D(k0b[13]),
    .Q(out_1[109]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _342_ (
    .C(clk),
    .CE(1'h1),
    .D(k0b[14]),
    .Q(out_1[110]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _343_ (
    .C(clk),
    .CE(1'h1),
    .D(k0b[15]),
    .Q(out_1[111]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _344_ (
    .C(clk),
    .CE(1'h1),
    .D(k0b[16]),
    .Q(out_1[112]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _345_ (
    .C(clk),
    .CE(1'h1),
    .D(k0b[17]),
    .Q(out_1[113]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _346_ (
    .C(clk),
    .CE(1'h1),
    .D(k0b[18]),
    .Q(out_1[114]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _347_ (
    .C(clk),
    .CE(1'h1),
    .D(k0b[19]),
    .Q(out_1[115]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _348_ (
    .C(clk),
    .CE(1'h1),
    .D(k0b[20]),
    .Q(out_1[116]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _349_ (
    .C(clk),
    .CE(1'h1),
    .D(k0b[21]),
    .Q(out_1[117]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _350_ (
    .C(clk),
    .CE(1'h1),
    .D(k0b[22]),
    .Q(out_1[118]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _351_ (
    .C(clk),
    .CE(1'h1),
    .D(k0b[23]),
    .Q(out_1[119]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _352_ (
    .C(clk),
    .CE(1'h1),
    .D(k0b[24]),
    .Q(out_1[120]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _353_ (
    .C(clk),
    .CE(1'h1),
    .D(k0b[25]),
    .Q(out_1[121]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _354_ (
    .C(clk),
    .CE(1'h1),
    .D(k0b[26]),
    .Q(out_1[122]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _355_ (
    .C(clk),
    .CE(1'h1),
    .D(k0b[27]),
    .Q(out_1[123]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _356_ (
    .C(clk),
    .CE(1'h1),
    .D(k0b[28]),
    .Q(out_1[124]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _357_ (
    .C(clk),
    .CE(1'h1),
    .D(k0b[29]),
    .Q(out_1[125]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _358_ (
    .C(clk),
    .CE(1'h1),
    .D(k0b[30]),
    .Q(out_1[126]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _359_ (
    .C(clk),
    .CE(1'h1),
    .D(k0b[31]),
    .Q(out_1[127]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _360_ (
    .C(clk),
    .CE(1'h1),
    .D(in[96]),
    .Q(k0a[0]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _361_ (
    .C(clk),
    .CE(1'h1),
    .D(in[97]),
    .Q(k0a[1]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _362_ (
    .C(clk),
    .CE(1'h1),
    .D(in[98]),
    .Q(k0a[2]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _363_ (
    .C(clk),
    .CE(1'h1),
    .D(in[99]),
    .Q(k0a[3]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _364_ (
    .C(clk),
    .CE(1'h1),
    .D(in[100]),
    .Q(k0a[4]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _365_ (
    .C(clk),
    .CE(1'h1),
    .D(in[101]),
    .Q(k0a[5]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _366_ (
    .C(clk),
    .CE(1'h1),
    .D(in[102]),
    .Q(k0a[6]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _367_ (
    .C(clk),
    .CE(1'h1),
    .D(in[103]),
    .Q(k0a[7]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _368_ (
    .C(clk),
    .CE(1'h1),
    .D(in[104]),
    .Q(k0a[8]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _369_ (
    .C(clk),
    .CE(1'h1),
    .D(in[105]),
    .Q(k0a[9]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _370_ (
    .C(clk),
    .CE(1'h1),
    .D(in[106]),
    .Q(k0a[10]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _371_ (
    .C(clk),
    .CE(1'h1),
    .D(in[107]),
    .Q(k0a[11]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _372_ (
    .C(clk),
    .CE(1'h1),
    .D(in[108]),
    .Q(k0a[12]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _373_ (
    .C(clk),
    .CE(1'h1),
    .D(in[109]),
    .Q(k0a[13]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _374_ (
    .C(clk),
    .CE(1'h1),
    .D(in[110]),
    .Q(k0a[14]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _375_ (
    .C(clk),
    .CE(1'h1),
    .D(in[111]),
    .Q(k0a[15]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _376_ (
    .C(clk),
    .CE(1'h1),
    .D(in[112]),
    .Q(k0a[16]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _377_ (
    .C(clk),
    .CE(1'h1),
    .D(in[113]),
    .Q(k0a[17]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _378_ (
    .C(clk),
    .CE(1'h1),
    .D(in[114]),
    .Q(k0a[18]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _379_ (
    .C(clk),
    .CE(1'h1),
    .D(in[115]),
    .Q(k0a[19]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _380_ (
    .C(clk),
    .CE(1'h1),
    .D(in[116]),
    .Q(k0a[20]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _381_ (
    .C(clk),
    .CE(1'h1),
    .D(in[117]),
    .Q(k0a[21]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _382_ (
    .C(clk),
    .CE(1'h1),
    .D(in[118]),
    .Q(k0a[22]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _383_ (
    .C(clk),
    .CE(1'h1),
    .D(in[119]),
    .Q(k0a[23]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _384_ (
    .C(clk),
    .CE(1'h1),
    .D(v0[24]),
    .Q(k0a[24]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _385_ (
    .C(clk),
    .CE(1'h1),
    .D(v0[25]),
    .Q(k0a[25]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _386_ (
    .C(clk),
    .CE(1'h1),
    .D(v0[26]),
    .Q(k0a[26]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _387_ (
    .C(clk),
    .CE(1'h1),
    .D(v0[27]),
    .Q(k0a[27]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _388_ (
    .C(clk),
    .CE(1'h1),
    .D(v0[28]),
    .Q(k0a[28]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _389_ (
    .C(clk),
    .CE(1'h1),
    .D(v0[29]),
    .Q(k0a[29]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _390_ (
    .C(clk),
    .CE(1'h1),
    .D(v0[30]),
    .Q(k0a[30]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _391_ (
    .C(clk),
    .CE(1'h1),
    .D(v0[31]),
    .Q(k0a[31]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _392_ (
    .C(clk),
    .CE(1'h1),
    .D(v1[0]),
    .Q(k1a[0]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _393_ (
    .C(clk),
    .CE(1'h1),
    .D(v1[1]),
    .Q(k1a[1]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _394_ (
    .C(clk),
    .CE(1'h1),
    .D(v1[2]),
    .Q(k1a[2]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _395_ (
    .C(clk),
    .CE(1'h1),
    .D(v1[3]),
    .Q(k1a[3]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _396_ (
    .C(clk),
    .CE(1'h1),
    .D(v1[4]),
    .Q(k1a[4]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _397_ (
    .C(clk),
    .CE(1'h1),
    .D(v1[5]),
    .Q(k1a[5]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _398_ (
    .C(clk),
    .CE(1'h1),
    .D(v1[6]),
    .Q(k1a[6]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _399_ (
    .C(clk),
    .CE(1'h1),
    .D(v1[7]),
    .Q(k1a[7]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _400_ (
    .C(clk),
    .CE(1'h1),
    .D(v1[8]),
    .Q(k1a[8]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _401_ (
    .C(clk),
    .CE(1'h1),
    .D(v1[9]),
    .Q(k1a[9]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _402_ (
    .C(clk),
    .CE(1'h1),
    .D(v1[10]),
    .Q(k1a[10]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _403_ (
    .C(clk),
    .CE(1'h1),
    .D(v1[11]),
    .Q(k1a[11]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _404_ (
    .C(clk),
    .CE(1'h1),
    .D(v1[12]),
    .Q(k1a[12]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _405_ (
    .C(clk),
    .CE(1'h1),
    .D(v1[13]),
    .Q(k1a[13]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _406_ (
    .C(clk),
    .CE(1'h1),
    .D(v1[14]),
    .Q(k1a[14]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _407_ (
    .C(clk),
    .CE(1'h1),
    .D(v1[15]),
    .Q(k1a[15]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _408_ (
    .C(clk),
    .CE(1'h1),
    .D(v1[16]),
    .Q(k1a[16]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _409_ (
    .C(clk),
    .CE(1'h1),
    .D(v1[17]),
    .Q(k1a[17]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _410_ (
    .C(clk),
    .CE(1'h1),
    .D(v1[18]),
    .Q(k1a[18]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _411_ (
    .C(clk),
    .CE(1'h1),
    .D(v1[19]),
    .Q(k1a[19]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _412_ (
    .C(clk),
    .CE(1'h1),
    .D(v1[20]),
    .Q(k1a[20]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _413_ (
    .C(clk),
    .CE(1'h1),
    .D(v1[21]),
    .Q(k1a[21]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _414_ (
    .C(clk),
    .CE(1'h1),
    .D(v1[22]),
    .Q(k1a[22]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _415_ (
    .C(clk),
    .CE(1'h1),
    .D(v1[23]),
    .Q(k1a[23]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _416_ (
    .C(clk),
    .CE(1'h1),
    .D(v1[24]),
    .Q(k1a[24]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _417_ (
    .C(clk),
    .CE(1'h1),
    .D(v1[25]),
    .Q(k1a[25]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _418_ (
    .C(clk),
    .CE(1'h1),
    .D(v1[26]),
    .Q(k1a[26]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _419_ (
    .C(clk),
    .CE(1'h1),
    .D(v1[27]),
    .Q(k1a[27]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _420_ (
    .C(clk),
    .CE(1'h1),
    .D(v1[28]),
    .Q(k1a[28]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _421_ (
    .C(clk),
    .CE(1'h1),
    .D(v1[29]),
    .Q(k1a[29]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _422_ (
    .C(clk),
    .CE(1'h1),
    .D(v1[30]),
    .Q(k1a[30]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _423_ (
    .C(clk),
    .CE(1'h1),
    .D(v1[31]),
    .Q(k1a[31]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _424_ (
    .C(clk),
    .CE(1'h1),
    .D(v2[0]),
    .Q(k2a[0]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _425_ (
    .C(clk),
    .CE(1'h1),
    .D(v2[1]),
    .Q(k2a[1]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _426_ (
    .C(clk),
    .CE(1'h1),
    .D(v2[2]),
    .Q(k2a[2]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _427_ (
    .C(clk),
    .CE(1'h1),
    .D(v2[3]),
    .Q(k2a[3]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _428_ (
    .C(clk),
    .CE(1'h1),
    .D(v2[4]),
    .Q(k2a[4]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _429_ (
    .C(clk),
    .CE(1'h1),
    .D(v2[5]),
    .Q(k2a[5]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _430_ (
    .C(clk),
    .CE(1'h1),
    .D(v2[6]),
    .Q(k2a[6]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _431_ (
    .C(clk),
    .CE(1'h1),
    .D(v2[7]),
    .Q(k2a[7]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _432_ (
    .C(clk),
    .CE(1'h1),
    .D(v2[8]),
    .Q(k2a[8]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _433_ (
    .C(clk),
    .CE(1'h1),
    .D(v2[9]),
    .Q(k2a[9]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _434_ (
    .C(clk),
    .CE(1'h1),
    .D(v2[10]),
    .Q(k2a[10]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _435_ (
    .C(clk),
    .CE(1'h1),
    .D(v2[11]),
    .Q(k2a[11]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _436_ (
    .C(clk),
    .CE(1'h1),
    .D(v2[12]),
    .Q(k2a[12]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _437_ (
    .C(clk),
    .CE(1'h1),
    .D(v2[13]),
    .Q(k2a[13]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _438_ (
    .C(clk),
    .CE(1'h1),
    .D(v2[14]),
    .Q(k2a[14]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _439_ (
    .C(clk),
    .CE(1'h1),
    .D(v2[15]),
    .Q(k2a[15]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _440_ (
    .C(clk),
    .CE(1'h1),
    .D(v2[16]),
    .Q(k2a[16]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _441_ (
    .C(clk),
    .CE(1'h1),
    .D(v2[17]),
    .Q(k2a[17]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _442_ (
    .C(clk),
    .CE(1'h1),
    .D(v2[18]),
    .Q(k2a[18]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _443_ (
    .C(clk),
    .CE(1'h1),
    .D(v2[19]),
    .Q(k2a[19]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _444_ (
    .C(clk),
    .CE(1'h1),
    .D(v2[20]),
    .Q(k2a[20]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _445_ (
    .C(clk),
    .CE(1'h1),
    .D(v2[21]),
    .Q(k2a[21]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _446_ (
    .C(clk),
    .CE(1'h1),
    .D(v2[22]),
    .Q(k2a[22]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _447_ (
    .C(clk),
    .CE(1'h1),
    .D(v2[23]),
    .Q(k2a[23]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _448_ (
    .C(clk),
    .CE(1'h1),
    .D(v2[24]),
    .Q(k2a[24]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _449_ (
    .C(clk),
    .CE(1'h1),
    .D(v2[25]),
    .Q(k2a[25]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _450_ (
    .C(clk),
    .CE(1'h1),
    .D(v2[26]),
    .Q(k2a[26]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _451_ (
    .C(clk),
    .CE(1'h1),
    .D(v2[27]),
    .Q(k2a[27]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _452_ (
    .C(clk),
    .CE(1'h1),
    .D(v2[28]),
    .Q(k2a[28]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _453_ (
    .C(clk),
    .CE(1'h1),
    .D(v2[29]),
    .Q(k2a[29]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _454_ (
    .C(clk),
    .CE(1'h1),
    .D(v2[30]),
    .Q(k2a[30]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _455_ (
    .C(clk),
    .CE(1'h1),
    .D(v2[31]),
    .Q(k2a[31]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _456_ (
    .C(clk),
    .CE(1'h1),
    .D(v3[0]),
    .Q(k3a[0]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _457_ (
    .C(clk),
    .CE(1'h1),
    .D(v3[1]),
    .Q(k3a[1]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _458_ (
    .C(clk),
    .CE(1'h1),
    .D(v3[2]),
    .Q(k3a[2]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _459_ (
    .C(clk),
    .CE(1'h1),
    .D(v3[3]),
    .Q(k3a[3]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _460_ (
    .C(clk),
    .CE(1'h1),
    .D(v3[4]),
    .Q(k3a[4]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _461_ (
    .C(clk),
    .CE(1'h1),
    .D(v3[5]),
    .Q(k3a[5]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _462_ (
    .C(clk),
    .CE(1'h1),
    .D(v3[6]),
    .Q(k3a[6]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _463_ (
    .C(clk),
    .CE(1'h1),
    .D(v3[7]),
    .Q(k3a[7]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _464_ (
    .C(clk),
    .CE(1'h1),
    .D(v3[8]),
    .Q(k3a[8]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _465_ (
    .C(clk),
    .CE(1'h1),
    .D(v3[9]),
    .Q(k3a[9]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _466_ (
    .C(clk),
    .CE(1'h1),
    .D(v3[10]),
    .Q(k3a[10]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _467_ (
    .C(clk),
    .CE(1'h1),
    .D(v3[11]),
    .Q(k3a[11]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _468_ (
    .C(clk),
    .CE(1'h1),
    .D(v3[12]),
    .Q(k3a[12]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _469_ (
    .C(clk),
    .CE(1'h1),
    .D(v3[13]),
    .Q(k3a[13]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _470_ (
    .C(clk),
    .CE(1'h1),
    .D(v3[14]),
    .Q(k3a[14]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _471_ (
    .C(clk),
    .CE(1'h1),
    .D(v3[15]),
    .Q(k3a[15]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _472_ (
    .C(clk),
    .CE(1'h1),
    .D(v3[16]),
    .Q(k3a[16]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _473_ (
    .C(clk),
    .CE(1'h1),
    .D(v3[17]),
    .Q(k3a[17]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _474_ (
    .C(clk),
    .CE(1'h1),
    .D(v3[18]),
    .Q(k3a[18]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _475_ (
    .C(clk),
    .CE(1'h1),
    .D(v3[19]),
    .Q(k3a[19]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _476_ (
    .C(clk),
    .CE(1'h1),
    .D(v3[20]),
    .Q(k3a[20]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _477_ (
    .C(clk),
    .CE(1'h1),
    .D(v3[21]),
    .Q(k3a[21]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _478_ (
    .C(clk),
    .CE(1'h1),
    .D(v3[22]),
    .Q(k3a[22]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _479_ (
    .C(clk),
    .CE(1'h1),
    .D(v3[23]),
    .Q(k3a[23]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _480_ (
    .C(clk),
    .CE(1'h1),
    .D(v3[24]),
    .Q(k3a[24]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _481_ (
    .C(clk),
    .CE(1'h1),
    .D(v3[25]),
    .Q(k3a[25]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _482_ (
    .C(clk),
    .CE(1'h1),
    .D(v3[26]),
    .Q(k3a[26]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _483_ (
    .C(clk),
    .CE(1'h1),
    .D(v3[27]),
    .Q(k3a[27]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _484_ (
    .C(clk),
    .CE(1'h1),
    .D(v3[28]),
    .Q(k3a[28]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _485_ (
    .C(clk),
    .CE(1'h1),
    .D(v3[29]),
    .Q(k3a[29]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _486_ (
    .C(clk),
    .CE(1'h1),
    .D(v3[30]),
    .Q(k3a[30]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _487_ (
    .C(clk),
    .CE(1'h1),
    .D(v3[31]),
    .Q(k3a[31]),
    .R(1'h0)
  );
S4  S4_0 (
    .clk(clk),
    .in({ in[23:0], in[31:24] }),
    .out(k4a)
  );
assign  k0 = in[127:96];
assign  k1 = in[95:64];
assign  k2 = in[63:32];
assign  k3 = in[31:0];
assign  out_2 = { k0b, k1b, k2b, k3b };
assign  v0[23:0] = in[119:96];
endmodule
