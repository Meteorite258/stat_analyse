module AES_Comp_EncCore(di,  ki, Rrg, \do , ko);
wire  [6:0] _000_;
wire  _001_;
wire  _002_;
wire  _003_;
wire  _004_;
wire  _005_;
wire  _006_;
wire  _007_;
wire  _008_;
wire  _009_;
wire  [6:0] _010_;
wire  _011_;
wire  _012_;
wire  _013_;
wire  _014_;
wire  _015_;
wire  _016_;
wire  _017_;
wire  _018_;
wire  _019_;
wire  [6:0] _020_;
wire  _021_;
wire  _022_;
wire  [6:0] _023_;
wire  _024_;
wire  _025_;
wire  [6:0] _026_;
wire  _027_;
wire  _028_;
wire  _029_;
wire  _030_;
wire  _031_;
wire  _032_;
wire  _033_;
wire  _034_;
wire  [6:0] _035_;
wire  _036_;
wire  _037_;
wire  [6:0] _038_;
wire  _039_;
wire  _040_;
wire  [6:0] _041_;
wire  _042_;
wire  _043_;
input  [9:0] Rrg;
wire  [9:0] Rrg;
input  [127:0] di;
wire  [127:0] di;
output  [127:0] \do ;
wire  [127:0] \do ;
input  [127:0] ki;
wire  [127:0] ki;
output  [127:0] ko;
wire  [127:0] ko;
wire  [127:0] mx;
wire  [9:0] \rcon$func$AES_Comp.v:349$425.x ;
wire  [127:0] sb;
wire  [31:0] so;
wire  [127:0] sr;
LUT4  #(
    .INIT(16'h53ac)
  ) _044_ (
    .I0(sb[9]),
    .I1(mx[73]),
    .I2(Rrg[0]),
    .I3(ki[73]),
    .O(\do [73])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _045_ (
    .I0(sb[10]),
    .I1(mx[74]),
    .I2(Rrg[0]),
    .I3(ki[74]),
    .O(\do [74])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _046_ (
    .I0(sb[11]),
    .I1(mx[75]),
    .I2(Rrg[0]),
    .I3(ki[75]),
    .O(\do [75])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _047_ (
    .I0(sb[12]),
    .I1(mx[76]),
    .I2(Rrg[0]),
    .I3(ki[76]),
    .O(\do [76])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _048_ (
    .I0(sb[13]),
    .I1(mx[77]),
    .I2(Rrg[0]),
    .I3(ki[77]),
    .O(\do [77])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _049_ (
    .I0(sb[14]),
    .I1(mx[78]),
    .I2(Rrg[0]),
    .I3(ki[78]),
    .O(\do [78])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _050_ (
    .I0(sb[15]),
    .I1(mx[79]),
    .I2(Rrg[0]),
    .I3(ki[79]),
    .O(\do [79])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _051_ (
    .I0(sb[48]),
    .I1(mx[80]),
    .I2(Rrg[0]),
    .I3(ki[80]),
    .O(\do [80])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _052_ (
    .I0(sb[49]),
    .I1(mx[81]),
    .I2(Rrg[0]),
    .I3(ki[81]),
    .O(\do [81])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _053_ (
    .I0(sb[50]),
    .I1(mx[82]),
    .I2(Rrg[0]),
    .I3(ki[82]),
    .O(\do [82])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _054_ (
    .I0(sb[51]),
    .I1(mx[83]),
    .I2(Rrg[0]),
    .I3(ki[83]),
    .O(\do [83])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _055_ (
    .I0(sb[52]),
    .I1(mx[84]),
    .I2(Rrg[0]),
    .I3(ki[84]),
    .O(\do [84])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _056_ (
    .I0(sb[53]),
    .I1(mx[85]),
    .I2(Rrg[0]),
    .I3(ki[85]),
    .O(\do [85])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _057_ (
    .I0(sb[54]),
    .I1(mx[86]),
    .I2(Rrg[0]),
    .I3(ki[86]),
    .O(\do [86])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _058_ (
    .I0(sb[55]),
    .I1(mx[87]),
    .I2(Rrg[0]),
    .I3(ki[87]),
    .O(\do [87])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _059_ (
    .I0(sb[88]),
    .I1(mx[88]),
    .I2(Rrg[0]),
    .I3(ki[88]),
    .O(\do [88])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _060_ (
    .I0(sb[89]),
    .I1(mx[89]),
    .I2(Rrg[0]),
    .I3(ki[89]),
    .O(\do [89])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _061_ (
    .I0(sb[90]),
    .I1(mx[90]),
    .I2(Rrg[0]),
    .I3(ki[90]),
    .O(\do [90])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _062_ (
    .I0(sb[91]),
    .I1(mx[91]),
    .I2(Rrg[0]),
    .I3(ki[91]),
    .O(\do [91])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _063_ (
    .I0(sb[92]),
    .I1(mx[92]),
    .I2(Rrg[0]),
    .I3(ki[92]),
    .O(\do [92])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _064_ (
    .I0(sb[93]),
    .I1(mx[93]),
    .I2(Rrg[0]),
    .I3(ki[93]),
    .O(\do [93])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _065_ (
    .I0(sb[94]),
    .I1(mx[94]),
    .I2(Rrg[0]),
    .I3(ki[94]),
    .O(\do [94])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _066_ (
    .I0(sb[95]),
    .I1(mx[95]),
    .I2(Rrg[0]),
    .I3(ki[95]),
    .O(\do [95])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _067_ (
    .I0(sb[0]),
    .I1(mx[96]),
    .I2(Rrg[0]),
    .I3(ki[96]),
    .O(\do [96])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _068_ (
    .I0(sb[1]),
    .I1(mx[97]),
    .I2(Rrg[0]),
    .I3(ki[97]),
    .O(\do [97])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _069_ (
    .I0(sb[2]),
    .I1(mx[98]),
    .I2(Rrg[0]),
    .I3(ki[98]),
    .O(\do [98])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _070_ (
    .I0(sb[3]),
    .I1(mx[99]),
    .I2(Rrg[0]),
    .I3(ki[99]),
    .O(\do [99])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _071_ (
    .I0(sb[4]),
    .I1(mx[100]),
    .I2(Rrg[0]),
    .I3(ki[100]),
    .O(\do [100])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _072_ (
    .I0(sb[5]),
    .I1(mx[101]),
    .I2(Rrg[0]),
    .I3(ki[101]),
    .O(\do [101])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _073_ (
    .I0(sb[6]),
    .I1(mx[102]),
    .I2(Rrg[0]),
    .I3(ki[102]),
    .O(\do [102])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _074_ (
    .I0(sb[7]),
    .I1(mx[103]),
    .I2(Rrg[0]),
    .I3(ki[103]),
    .O(\do [103])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _075_ (
    .I0(sb[40]),
    .I1(mx[104]),
    .I2(Rrg[0]),
    .I3(ki[104]),
    .O(\do [104])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _076_ (
    .I0(sb[41]),
    .I1(mx[105]),
    .I2(Rrg[0]),
    .I3(ki[105]),
    .O(\do [105])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _077_ (
    .I0(sb[42]),
    .I1(mx[106]),
    .I2(Rrg[0]),
    .I3(ki[106]),
    .O(\do [106])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _078_ (
    .I0(sb[43]),
    .I1(mx[107]),
    .I2(Rrg[0]),
    .I3(ki[107]),
    .O(\do [107])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _079_ (
    .I0(sb[44]),
    .I1(mx[108]),
    .I2(Rrg[0]),
    .I3(ki[108]),
    .O(\do [108])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _080_ (
    .I0(sb[45]),
    .I1(mx[109]),
    .I2(Rrg[0]),
    .I3(ki[109]),
    .O(\do [109])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _081_ (
    .I0(sb[46]),
    .I1(mx[110]),
    .I2(Rrg[0]),
    .I3(ki[110]),
    .O(\do [110])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _082_ (
    .I0(sb[47]),
    .I1(mx[111]),
    .I2(Rrg[0]),
    .I3(ki[111]),
    .O(\do [111])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _083_ (
    .I0(sb[80]),
    .I1(mx[112]),
    .I2(Rrg[0]),
    .I3(ki[112]),
    .O(\do [112])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _084_ (
    .I0(sb[81]),
    .I1(mx[113]),
    .I2(Rrg[0]),
    .I3(ki[113]),
    .O(\do [113])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _085_ (
    .I0(sb[82]),
    .I1(mx[114]),
    .I2(Rrg[0]),
    .I3(ki[114]),
    .O(\do [114])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _086_ (
    .I0(sb[83]),
    .I1(mx[115]),
    .I2(Rrg[0]),
    .I3(ki[115]),
    .O(\do [115])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _087_ (
    .I0(sb[84]),
    .I1(mx[116]),
    .I2(Rrg[0]),
    .I3(ki[116]),
    .O(\do [116])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _088_ (
    .I0(sb[85]),
    .I1(mx[117]),
    .I2(Rrg[0]),
    .I3(ki[117]),
    .O(\do [117])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _089_ (
    .I0(sb[86]),
    .I1(mx[118]),
    .I2(Rrg[0]),
    .I3(ki[118]),
    .O(\do [118])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _090_ (
    .I0(sb[87]),
    .I1(mx[119]),
    .I2(Rrg[0]),
    .I3(ki[119]),
    .O(\do [119])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _091_ (
    .I0(sb[120]),
    .I1(mx[120]),
    .I2(Rrg[0]),
    .I3(ki[120]),
    .O(\do [120])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _092_ (
    .I0(sb[121]),
    .I1(mx[121]),
    .I2(Rrg[0]),
    .I3(ki[121]),
    .O(\do [121])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _093_ (
    .I0(sb[122]),
    .I1(mx[122]),
    .I2(Rrg[0]),
    .I3(ki[122]),
    .O(\do [122])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _094_ (
    .I0(sb[123]),
    .I1(mx[123]),
    .I2(Rrg[0]),
    .I3(ki[123]),
    .O(\do [123])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _095_ (
    .I0(sb[124]),
    .I1(mx[124]),
    .I2(Rrg[0]),
    .I3(ki[124]),
    .O(\do [124])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _096_ (
    .I0(sb[125]),
    .I1(mx[125]),
    .I2(Rrg[0]),
    .I3(ki[125]),
    .O(\do [125])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _097_ (
    .I0(sb[126]),
    .I1(mx[126]),
    .I2(Rrg[0]),
    .I3(ki[126]),
    .O(\do [126])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _098_ (
    .I0(sb[127]),
    .I1(mx[127]),
    .I2(Rrg[0]),
    .I3(ki[127]),
    .O(\do [127])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _099_ (
    .I0(ki[32]),
    .I1(ki[64]),
    .I2(ki[96]),
    .I3(so[0]),
    .O(ko[32])
  );
LUT2  #(
    .INIT(4'h6)
  ) _100_ (
    .I0(ko[32]),
    .I1(ki[0]),
    .O(ko[0])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _101_ (
    .I0(ki[33]),
    .I1(ki[65]),
    .I2(ki[97]),
    .I3(so[1]),
    .O(ko[33])
  );
LUT2  #(
    .INIT(4'h6)
  ) _102_ (
    .I0(ko[33]),
    .I1(ki[1]),
    .O(ko[1])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _103_ (
    .I0(ki[34]),
    .I1(ki[66]),
    .I2(ki[98]),
    .I3(so[2]),
    .O(ko[34])
  );
LUT2  #(
    .INIT(4'h6)
  ) _104_ (
    .I0(ko[34]),
    .I1(ki[2]),
    .O(ko[2])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _105_ (
    .I0(ki[35]),
    .I1(ki[67]),
    .I2(ki[99]),
    .I3(so[3]),
    .O(ko[35])
  );
LUT2  #(
    .INIT(4'h6)
  ) _106_ (
    .I0(ko[35]),
    .I1(ki[3]),
    .O(ko[3])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _107_ (
    .I0(ki[36]),
    .I1(ki[68]),
    .I2(ki[100]),
    .I3(so[4]),
    .O(ko[36])
  );
LUT2  #(
    .INIT(4'h6)
  ) _108_ (
    .I0(ko[36]),
    .I1(ki[4]),
    .O(ko[4])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _109_ (
    .I0(ki[37]),
    .I1(ki[69]),
    .I2(ki[101]),
    .I3(so[5]),
    .O(ko[37])
  );
LUT2  #(
    .INIT(4'h6)
  ) _110_ (
    .I0(ko[37]),
    .I1(ki[5]),
    .O(ko[5])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _111_ (
    .I0(ki[38]),
    .I1(ki[70]),
    .I2(ki[102]),
    .I3(so[6]),
    .O(ko[38])
  );
LUT2  #(
    .INIT(4'h6)
  ) _112_ (
    .I0(ko[38]),
    .I1(ki[6]),
    .O(ko[6])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _113_ (
    .I0(ki[39]),
    .I1(ki[71]),
    .I2(ki[103]),
    .I3(so[7]),
    .O(ko[39])
  );
LUT2  #(
    .INIT(4'h6)
  ) _114_ (
    .I0(ko[39]),
    .I1(ki[7]),
    .O(ko[7])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _115_ (
    .I0(ki[40]),
    .I1(ki[72]),
    .I2(ki[104]),
    .I3(so[8]),
    .O(ko[40])
  );
LUT2  #(
    .INIT(4'h6)
  ) _116_ (
    .I0(ko[40]),
    .I1(ki[8]),
    .O(ko[8])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _117_ (
    .I0(ki[41]),
    .I1(ki[73]),
    .I2(ki[105]),
    .I3(so[9]),
    .O(ko[41])
  );
LUT2  #(
    .INIT(4'h6)
  ) _118_ (
    .I0(ko[41]),
    .I1(ki[9]),
    .O(ko[9])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _119_ (
    .I0(ki[42]),
    .I1(ki[74]),
    .I2(ki[106]),
    .I3(so[10]),
    .O(ko[42])
  );
LUT2  #(
    .INIT(4'h6)
  ) _120_ (
    .I0(ko[42]),
    .I1(ki[10]),
    .O(ko[10])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _121_ (
    .I0(ki[43]),
    .I1(ki[75]),
    .I2(ki[107]),
    .I3(so[11]),
    .O(ko[43])
  );
LUT2  #(
    .INIT(4'h6)
  ) _122_ (
    .I0(ko[43]),
    .I1(ki[11]),
    .O(ko[11])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _123_ (
    .I0(ki[44]),
    .I1(ki[76]),
    .I2(ki[108]),
    .I3(so[12]),
    .O(ko[44])
  );
LUT2  #(
    .INIT(4'h6)
  ) _124_ (
    .I0(ko[44]),
    .I1(ki[12]),
    .O(ko[12])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _125_ (
    .I0(ki[45]),
    .I1(ki[77]),
    .I2(ki[109]),
    .I3(so[13]),
    .O(ko[45])
  );
LUT2  #(
    .INIT(4'h6)
  ) _126_ (
    .I0(ko[45]),
    .I1(ki[13]),
    .O(ko[13])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _127_ (
    .I0(ki[46]),
    .I1(ki[78]),
    .I2(ki[110]),
    .I3(so[14]),
    .O(ko[46])
  );
LUT2  #(
    .INIT(4'h6)
  ) _128_ (
    .I0(ko[46]),
    .I1(ki[14]),
    .O(ko[14])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _129_ (
    .I0(ki[47]),
    .I1(ki[79]),
    .I2(ki[111]),
    .I3(so[15]),
    .O(ko[47])
  );
LUT2  #(
    .INIT(4'h6)
  ) _130_ (
    .I0(ko[47]),
    .I1(ki[15]),
    .O(ko[15])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _131_ (
    .I0(ki[48]),
    .I1(ki[80]),
    .I2(ki[112]),
    .I3(so[16]),
    .O(ko[48])
  );
LUT2  #(
    .INIT(4'h6)
  ) _132_ (
    .I0(ko[48]),
    .I1(ki[16]),
    .O(ko[16])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _133_ (
    .I0(ki[49]),
    .I1(ki[81]),
    .I2(ki[113]),
    .I3(so[17]),
    .O(ko[49])
  );
LUT2  #(
    .INIT(4'h6)
  ) _134_ (
    .I0(ko[49]),
    .I1(ki[17]),
    .O(ko[17])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _135_ (
    .I0(ki[50]),
    .I1(ki[82]),
    .I2(ki[114]),
    .I3(so[18]),
    .O(ko[50])
  );
LUT2  #(
    .INIT(4'h6)
  ) _136_ (
    .I0(ko[50]),
    .I1(ki[18]),
    .O(ko[18])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _137_ (
    .I0(ki[51]),
    .I1(ki[83]),
    .I2(ki[115]),
    .I3(so[19]),
    .O(ko[51])
  );
LUT2  #(
    .INIT(4'h6)
  ) _138_ (
    .I0(ko[51]),
    .I1(ki[19]),
    .O(ko[19])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _139_ (
    .I0(ki[52]),
    .I1(ki[84]),
    .I2(ki[116]),
    .I3(so[20]),
    .O(ko[52])
  );
LUT2  #(
    .INIT(4'h6)
  ) _140_ (
    .I0(ko[52]),
    .I1(ki[20]),
    .O(ko[20])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _141_ (
    .I0(ki[53]),
    .I1(ki[85]),
    .I2(ki[117]),
    .I3(so[21]),
    .O(ko[53])
  );
LUT2  #(
    .INIT(4'h6)
  ) _142_ (
    .I0(ko[53]),
    .I1(ki[21]),
    .O(ko[21])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _143_ (
    .I0(ki[54]),
    .I1(ki[86]),
    .I2(ki[118]),
    .I3(so[22]),
    .O(ko[54])
  );
LUT2  #(
    .INIT(4'h6)
  ) _144_ (
    .I0(ko[54]),
    .I1(ki[22]),
    .O(ko[22])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _145_ (
    .I0(ki[55]),
    .I1(ki[87]),
    .I2(ki[119]),
    .I3(so[23]),
    .O(ko[55])
  );
LUT2  #(
    .INIT(4'h6)
  ) _146_ (
    .I0(ko[55]),
    .I1(ki[23]),
    .O(ko[23])
  );
LUT6  #(
    .INIT(64'h07f8f807f80707f8)
  ) _147_ (
    .I0(_000_[0]),
    .I1(Rrg[8]),
    .I2(Rrg[0]),
    .I3(ki[56]),
    .I4(ki[88]),
    .I5(ki[120]),
    .O(_001_)
  );
LUT6  #(
    .INIT(64'hf80707f807f8f807)
  ) _148_ (
    .I0(_000_[0]),
    .I1(Rrg[8]),
    .I2(Rrg[0]),
    .I3(ki[56]),
    .I4(ki[88]),
    .I5(ki[120]),
    .O(_002_)
  );
MUXF7  _149_ (
    .I0(_001_),
    .I1(_002_),
    .O(ko[56]),
    .S(so[24])
  );
LUT6  #(
    .INIT(64'h0000000000000001)
  ) _150_ (
    .I0(Rrg[7]),
    .I1(Rrg[6]),
    .I2(Rrg[5]),
    .I3(Rrg[4]),
    .I4(Rrg[3]),
    .I5(Rrg[2]),
    .O(_003_)
  );
MUXF7  _151_ (
    .I0(_003_),
    .I1(1'h0),
    .O(_000_[0]),
    .S(Rrg[1])
  );
LUT6  #(
    .INIT(64'h07f8f807f80707f8)
  ) _152_ (
    .I0(_000_[0]),
    .I1(Rrg[8]),
    .I2(Rrg[0]),
    .I3(ki[24]),
    .I4(ki[56]),
    .I5(ki[88]),
    .O(_006_)
  );
LUT6  #(
    .INIT(64'hf80707f807f8f807)
  ) _153_ (
    .I0(_000_[0]),
    .I1(Rrg[8]),
    .I2(Rrg[0]),
    .I3(ki[24]),
    .I4(ki[56]),
    .I5(ki[88]),
    .O(_007_)
  );
MUXF7  _154_ (
    .I0(_006_),
    .I1(_007_),
    .O(_004_),
    .S(ki[120])
  );
LUT6  #(
    .INIT(64'hf80707f807f8f807)
  ) _155_ (
    .I0(_000_[0]),
    .I1(Rrg[8]),
    .I2(Rrg[0]),
    .I3(ki[24]),
    .I4(ki[56]),
    .I5(ki[88]),
    .O(_008_)
  );
LUT6  #(
    .INIT(64'h07f8f807f80707f8)
  ) _156_ (
    .I0(_000_[0]),
    .I1(Rrg[8]),
    .I2(Rrg[0]),
    .I3(ki[24]),
    .I4(ki[56]),
    .I5(ki[88]),
    .O(_009_)
  );
MUXF7  _157_ (
    .I0(_008_),
    .I1(_009_),
    .O(_005_),
    .S(ki[120])
  );
MUXF8  _158_ (
    .I0(_004_),
    .I1(_005_),
    .O(ko[24]),
    .S(so[24])
  );
LUT6  #(
    .INIT(64'hf10e0ef10ef1f10e)
  ) _159_ (
    .I0(_010_[0]),
    .I1(Rrg[1]),
    .I2(Rrg[0]),
    .I3(ki[57]),
    .I4(ki[89]),
    .I5(ki[121]),
    .O(_011_)
  );
LUT6  #(
    .INIT(64'h0ef1f10ef10e0ef1)
  ) _160_ (
    .I0(_010_[0]),
    .I1(Rrg[1]),
    .I2(Rrg[0]),
    .I3(ki[57]),
    .I4(ki[89]),
    .I5(ki[121]),
    .O(_012_)
  );
MUXF7  _161_ (
    .I0(_011_),
    .I1(_012_),
    .O(ko[57]),
    .S(so[25])
  );
LUT6  #(
    .INIT(64'h0000000000000001)
  ) _162_ (
    .I0(Rrg[7]),
    .I1(Rrg[6]),
    .I2(Rrg[5]),
    .I3(Rrg[4]),
    .I4(Rrg[3]),
    .I5(Rrg[2]),
    .O(_010_[0])
  );
LUT6  #(
    .INIT(64'hf10e0ef10ef1f10e)
  ) _163_ (
    .I0(_010_[0]),
    .I1(Rrg[1]),
    .I2(Rrg[0]),
    .I3(ki[25]),
    .I4(ki[57]),
    .I5(ki[89]),
    .O(_015_)
  );
LUT6  #(
    .INIT(64'h0ef1f10ef10e0ef1)
  ) _164_ (
    .I0(_010_[0]),
    .I1(Rrg[1]),
    .I2(Rrg[0]),
    .I3(ki[25]),
    .I4(ki[57]),
    .I5(ki[89]),
    .O(_016_)
  );
MUXF7  _165_ (
    .I0(_015_),
    .I1(_016_),
    .O(_013_),
    .S(ki[121])
  );
LUT6  #(
    .INIT(64'h0ef1f10ef10e0ef1)
  ) _166_ (
    .I0(_010_[0]),
    .I1(Rrg[1]),
    .I2(Rrg[0]),
    .I3(ki[25]),
    .I4(ki[57]),
    .I5(ki[89]),
    .O(_017_)
  );
LUT6  #(
    .INIT(64'hf10e0ef10ef1f10e)
  ) _167_ (
    .I0(_010_[0]),
    .I1(Rrg[1]),
    .I2(Rrg[0]),
    .I3(ki[25]),
    .I4(ki[57]),
    .I5(ki[89]),
    .O(_018_)
  );
MUXF7  _168_ (
    .I0(_017_),
    .I1(_018_),
    .O(_014_),
    .S(ki[121])
  );
MUXF8  _169_ (
    .I0(_013_),
    .I1(_014_),
    .O(ko[25]),
    .S(so[25])
  );
LUT6  #(
    .INIT(64'h4bb4b44bb44b4bb4)
  ) _170_ (
    .I0(_020_[0]),
    .I1(_020_[1]),
    .I2(ki[58]),
    .I3(ki[90]),
    .I4(ki[122]),
    .I5(so[26]),
    .O(ko[58])
  );
LUT6  #(
    .INIT(64'hfffffffffffffffe)
  ) _171_ (
    .I0(Rrg[7]),
    .I1(Rrg[6]),
    .I2(Rrg[5]),
    .I3(Rrg[4]),
    .I4(Rrg[3]),
    .I5(Rrg[8]),
    .O(_019_)
  );
MUXF7  _172_ (
    .I0(_019_),
    .I1(1'h0),
    .O(_020_[0]),
    .S(Rrg[2])
  );
LUT2  #(
    .INIT(4'h1)
  ) _173_ (
    .I0(Rrg[0]),
    .I1(Rrg[1]),
    .O(_020_[1])
  );
LUT6  #(
    .INIT(64'h4bb4b44bb44b4bb4)
  ) _174_ (
    .I0(_020_[0]),
    .I1(_020_[1]),
    .I2(ki[26]),
    .I3(ki[58]),
    .I4(ki[90]),
    .I5(ki[122]),
    .O(_021_)
  );
LUT6  #(
    .INIT(64'hb44b4bb44bb4b44b)
  ) _175_ (
    .I0(_020_[0]),
    .I1(_020_[1]),
    .I2(ki[26]),
    .I3(ki[58]),
    .I4(ki[90]),
    .I5(ki[122]),
    .O(_022_)
  );
MUXF7  _176_ (
    .I0(_021_),
    .I1(_022_),
    .O(ko[26]),
    .S(so[26])
  );
LUT6  #(
    .INIT(64'h4bb4b44bb44b4bb4)
  ) _177_ (
    .I0(_023_[0]),
    .I1(_023_[1]),
    .I2(ki[59]),
    .I3(ki[91]),
    .I4(ki[123]),
    .I5(so[27]),
    .O(ko[59])
  );
LUT6  #(
    .INIT(64'h00000000fffeffff)
  ) _178_ (
    .I0(Rrg[7]),
    .I1(Rrg[6]),
    .I2(Rrg[5]),
    .I3(Rrg[4]),
    .I4(Rrg[8]),
    .I5(Rrg[3]),
    .O(_023_[0])
  );
LUT3  #(
    .INIT(8'h01)
  ) _179_ (
    .I0(Rrg[0]),
    .I1(Rrg[2]),
    .I2(Rrg[1]),
    .O(_023_[1])
  );
LUT6  #(
    .INIT(64'h4bb4b44bb44b4bb4)
  ) _180_ (
    .I0(_023_[0]),
    .I1(_023_[1]),
    .I2(ki[27]),
    .I3(ki[59]),
    .I4(ki[91]),
    .I5(ki[123]),
    .O(_024_)
  );
LUT6  #(
    .INIT(64'hb44b4bb44bb4b44b)
  ) _181_ (
    .I0(_023_[0]),
    .I1(_023_[1]),
    .I2(ki[27]),
    .I3(ki[59]),
    .I4(ki[91]),
    .I5(ki[123]),
    .O(_025_)
  );
MUXF7  _182_ (
    .I0(_024_),
    .I1(_025_),
    .O(ko[27]),
    .S(so[27])
  );
LUT6  #(
    .INIT(64'h1fe0e01fe01f1fe0)
  ) _183_ (
    .I0(_026_[0]),
    .I1(Rrg[4]),
    .I2(_026_[2]),
    .I3(ki[60]),
    .I4(ki[92]),
    .I5(ki[124]),
    .O(_027_)
  );
LUT6  #(
    .INIT(64'he01f1fe01fe0e01f)
  ) _184_ (
    .I0(_026_[0]),
    .I1(Rrg[4]),
    .I2(_026_[2]),
    .I3(ki[60]),
    .I4(ki[92]),
    .I5(ki[124]),
    .O(_028_)
  );
MUXF7  _185_ (
    .I0(_027_),
    .I1(_028_),
    .O(ko[60]),
    .S(so[28])
  );
LUT3  #(
    .INIT(8'h01)
  ) _186_ (
    .I0(Rrg[7]),
    .I1(Rrg[6]),
    .I2(Rrg[5]),
    .O(_026_[0])
  );
LUT4  #(
    .INIT(16'h0001)
  ) _187_ (
    .I0(Rrg[0]),
    .I1(Rrg[3]),
    .I2(Rrg[2]),
    .I3(Rrg[1]),
    .O(_026_[2])
  );
LUT6  #(
    .INIT(64'h1fe0e01fe01f1fe0)
  ) _188_ (
    .I0(_026_[0]),
    .I1(Rrg[4]),
    .I2(_026_[2]),
    .I3(ki[28]),
    .I4(ki[60]),
    .I5(ki[92]),
    .O(_031_)
  );
LUT6  #(
    .INIT(64'he01f1fe01fe0e01f)
  ) _189_ (
    .I0(_026_[0]),
    .I1(Rrg[4]),
    .I2(_026_[2]),
    .I3(ki[28]),
    .I4(ki[60]),
    .I5(ki[92]),
    .O(_032_)
  );
MUXF7  _190_ (
    .I0(_031_),
    .I1(_032_),
    .O(_029_),
    .S(ki[124])
  );
LUT6  #(
    .INIT(64'he01f1fe01fe0e01f)
  ) _191_ (
    .I0(_026_[0]),
    .I1(Rrg[4]),
    .I2(_026_[2]),
    .I3(ki[28]),
    .I4(ki[60]),
    .I5(ki[92]),
    .O(_033_)
  );
LUT6  #(
    .INIT(64'h1fe0e01fe01f1fe0)
  ) _192_ (
    .I0(_026_[0]),
    .I1(Rrg[4]),
    .I2(_026_[2]),
    .I3(ki[28]),
    .I4(ki[60]),
    .I5(ki[92]),
    .O(_034_)
  );
MUXF7  _193_ (
    .I0(_033_),
    .I1(_034_),
    .O(_030_),
    .S(ki[124])
  );
MUXF8  _194_ (
    .I0(_029_),
    .I1(_030_),
    .O(ko[28]),
    .S(so[28])
  );
LUT6  #(
    .INIT(64'h4bb4b44bb44b4bb4)
  ) _195_ (
    .I0(_035_[0]),
    .I1(_035_[1]),
    .I2(ki[61]),
    .I3(ki[93]),
    .I4(ki[125]),
    .I5(so[29]),
    .O(ko[61])
  );
LUT4  #(
    .INIT(16'h00fe)
  ) _196_ (
    .I0(Rrg[7]),
    .I1(Rrg[6]),
    .I2(Rrg[8]),
    .I3(Rrg[5]),
    .O(_035_[0])
  );
LUT5  #(
    .INIT(32'd1)
  ) _197_ (
    .I0(Rrg[0]),
    .I1(Rrg[4]),
    .I2(Rrg[3]),
    .I3(Rrg[2]),
    .I4(Rrg[1]),
    .O(_035_[1])
  );
LUT6  #(
    .INIT(64'h4bb4b44bb44b4bb4)
  ) _198_ (
    .I0(_035_[0]),
    .I1(_035_[1]),
    .I2(ki[29]),
    .I3(ki[61]),
    .I4(ki[93]),
    .I5(ki[125]),
    .O(_036_)
  );
LUT6  #(
    .INIT(64'hb44b4bb44bb4b44b)
  ) _199_ (
    .I0(_035_[0]),
    .I1(_035_[1]),
    .I2(ki[29]),
    .I3(ki[61]),
    .I4(ki[93]),
    .I5(ki[125]),
    .O(_037_)
  );
MUXF7  _200_ (
    .I0(_036_),
    .I1(_037_),
    .O(ko[29]),
    .S(so[29])
  );
LUT6  #(
    .INIT(64'h8778788778878778)
  ) _201_ (
    .I0(_035_[1]),
    .I1(_038_[1]),
    .I2(ki[62]),
    .I3(ki[94]),
    .I4(ki[126]),
    .I5(so[30]),
    .O(ko[62])
  );
LUT2  #(
    .INIT(4'h4)
  ) _202_ (
    .I0(Rrg[5]),
    .I1(Rrg[6]),
    .O(_038_[1])
  );
LUT6  #(
    .INIT(64'h8778788778878778)
  ) _203_ (
    .I0(_035_[1]),
    .I1(_038_[1]),
    .I2(ki[30]),
    .I3(ki[62]),
    .I4(ki[94]),
    .I5(ki[126]),
    .O(_039_)
  );
LUT6  #(
    .INIT(64'h7887877887787887)
  ) _204_ (
    .I0(_035_[1]),
    .I1(_038_[1]),
    .I2(ki[30]),
    .I3(ki[62]),
    .I4(ki[94]),
    .I5(ki[126]),
    .O(_040_)
  );
MUXF7  _205_ (
    .I0(_039_),
    .I1(_040_),
    .O(ko[30]),
    .S(so[30])
  );
LUT6  #(
    .INIT(64'h8778788778878778)
  ) _206_ (
    .I0(_035_[1]),
    .I1(_041_[1]),
    .I2(ki[63]),
    .I3(ki[95]),
    .I4(ki[127]),
    .I5(so[31]),
    .O(ko[63])
  );
LUT3  #(
    .INIT(8'h10)
  ) _207_ (
    .I0(Rrg[6]),
    .I1(Rrg[5]),
    .I2(Rrg[7]),
    .O(_041_[1])
  );
LUT6  #(
    .INIT(64'h8778788778878778)
  ) _208_ (
    .I0(_035_[1]),
    .I1(_041_[1]),
    .I2(ki[31]),
    .I3(ki[63]),
    .I4(ki[95]),
    .I5(ki[127]),
    .O(_042_)
  );
LUT6  #(
    .INIT(64'h7887877887787887)
  ) _209_ (
    .I0(_035_[1]),
    .I1(_041_[1]),
    .I2(ki[31]),
    .I3(ki[63]),
    .I4(ki[95]),
    .I5(ki[127]),
    .O(_043_)
  );
MUXF7  _210_ (
    .I0(_042_),
    .I1(_043_),
    .O(ko[31]),
    .S(so[31])
  );
LUT2  #(
    .INIT(4'h6)
  ) _211_ (
    .I0(ko[96]),
    .I1(ki[64]),
    .O(ko[64])
  );
LUT2  #(
    .INIT(4'h6)
  ) _212_ (
    .I0(ki[96]),
    .I1(so[0]),
    .O(ko[96])
  );
LUT2  #(
    .INIT(4'h6)
  ) _213_ (
    .I0(ko[97]),
    .I1(ki[65]),
    .O(ko[65])
  );
LUT2  #(
    .INIT(4'h6)
  ) _214_ (
    .I0(ki[97]),
    .I1(so[1]),
    .O(ko[97])
  );
LUT2  #(
    .INIT(4'h6)
  ) _215_ (
    .I0(ko[98]),
    .I1(ki[66]),
    .O(ko[66])
  );
LUT2  #(
    .INIT(4'h6)
  ) _216_ (
    .I0(ki[98]),
    .I1(so[2]),
    .O(ko[98])
  );
LUT2  #(
    .INIT(4'h6)
  ) _217_ (
    .I0(ko[99]),
    .I1(ki[67]),
    .O(ko[67])
  );
LUT2  #(
    .INIT(4'h6)
  ) _218_ (
    .I0(ki[99]),
    .I1(so[3]),
    .O(ko[99])
  );
LUT2  #(
    .INIT(4'h6)
  ) _219_ (
    .I0(ko[100]),
    .I1(ki[68]),
    .O(ko[68])
  );
LUT2  #(
    .INIT(4'h6)
  ) _220_ (
    .I0(ki[100]),
    .I1(so[4]),
    .O(ko[100])
  );
LUT2  #(
    .INIT(4'h6)
  ) _221_ (
    .I0(ko[101]),
    .I1(ki[69]),
    .O(ko[69])
  );
LUT2  #(
    .INIT(4'h6)
  ) _222_ (
    .I0(ki[101]),
    .I1(so[5]),
    .O(ko[101])
  );
LUT2  #(
    .INIT(4'h6)
  ) _223_ (
    .I0(ko[102]),
    .I1(ki[70]),
    .O(ko[70])
  );
LUT2  #(
    .INIT(4'h6)
  ) _224_ (
    .I0(ki[102]),
    .I1(so[6]),
    .O(ko[102])
  );
LUT2  #(
    .INIT(4'h6)
  ) _225_ (
    .I0(ko[103]),
    .I1(ki[71]),
    .O(ko[71])
  );
LUT2  #(
    .INIT(4'h6)
  ) _226_ (
    .I0(ki[103]),
    .I1(so[7]),
    .O(ko[103])
  );
LUT2  #(
    .INIT(4'h6)
  ) _227_ (
    .I0(ko[104]),
    .I1(ki[72]),
    .O(ko[72])
  );
LUT2  #(
    .INIT(4'h6)
  ) _228_ (
    .I0(ki[104]),
    .I1(so[8]),
    .O(ko[104])
  );
LUT2  #(
    .INIT(4'h6)
  ) _229_ (
    .I0(ko[105]),
    .I1(ki[73]),
    .O(ko[73])
  );
LUT2  #(
    .INIT(4'h6)
  ) _230_ (
    .I0(ki[105]),
    .I1(so[9]),
    .O(ko[105])
  );
LUT2  #(
    .INIT(4'h6)
  ) _231_ (
    .I0(ko[106]),
    .I1(ki[74]),
    .O(ko[74])
  );
LUT2  #(
    .INIT(4'h6)
  ) _232_ (
    .I0(ki[106]),
    .I1(so[10]),
    .O(ko[106])
  );
LUT2  #(
    .INIT(4'h6)
  ) _233_ (
    .I0(ko[107]),
    .I1(ki[75]),
    .O(ko[75])
  );
LUT2  #(
    .INIT(4'h6)
  ) _234_ (
    .I0(ki[107]),
    .I1(so[11]),
    .O(ko[107])
  );
LUT2  #(
    .INIT(4'h6)
  ) _235_ (
    .I0(ko[108]),
    .I1(ki[76]),
    .O(ko[76])
  );
LUT2  #(
    .INIT(4'h6)
  ) _236_ (
    .I0(ki[108]),
    .I1(so[12]),
    .O(ko[108])
  );
LUT2  #(
    .INIT(4'h6)
  ) _237_ (
    .I0(ko[109]),
    .I1(ki[77]),
    .O(ko[77])
  );
LUT2  #(
    .INIT(4'h6)
  ) _238_ (
    .I0(ki[109]),
    .I1(so[13]),
    .O(ko[109])
  );
LUT2  #(
    .INIT(4'h6)
  ) _239_ (
    .I0(ko[110]),
    .I1(ki[78]),
    .O(ko[78])
  );
LUT2  #(
    .INIT(4'h6)
  ) _240_ (
    .I0(ki[110]),
    .I1(so[14]),
    .O(ko[110])
  );
LUT2  #(
    .INIT(4'h6)
  ) _241_ (
    .I0(ko[111]),
    .I1(ki[79]),
    .O(ko[79])
  );
LUT2  #(
    .INIT(4'h6)
  ) _242_ (
    .I0(ki[111]),
    .I1(so[15]),
    .O(ko[111])
  );
LUT2  #(
    .INIT(4'h6)
  ) _243_ (
    .I0(ko[112]),
    .I1(ki[80]),
    .O(ko[80])
  );
LUT2  #(
    .INIT(4'h6)
  ) _244_ (
    .I0(ki[112]),
    .I1(so[16]),
    .O(ko[112])
  );
LUT2  #(
    .INIT(4'h6)
  ) _245_ (
    .I0(ko[113]),
    .I1(ki[81]),
    .O(ko[81])
  );
LUT2  #(
    .INIT(4'h6)
  ) _246_ (
    .I0(ki[113]),
    .I1(so[17]),
    .O(ko[113])
  );
LUT2  #(
    .INIT(4'h6)
  ) _247_ (
    .I0(ko[114]),
    .I1(ki[82]),
    .O(ko[82])
  );
LUT2  #(
    .INIT(4'h6)
  ) _248_ (
    .I0(ki[114]),
    .I1(so[18]),
    .O(ko[114])
  );
LUT2  #(
    .INIT(4'h6)
  ) _249_ (
    .I0(ko[115]),
    .I1(ki[83]),
    .O(ko[83])
  );
LUT2  #(
    .INIT(4'h6)
  ) _250_ (
    .I0(ki[115]),
    .I1(so[19]),
    .O(ko[115])
  );
LUT2  #(
    .INIT(4'h6)
  ) _251_ (
    .I0(ko[116]),
    .I1(ki[84]),
    .O(ko[84])
  );
LUT2  #(
    .INIT(4'h6)
  ) _252_ (
    .I0(ki[116]),
    .I1(so[20]),
    .O(ko[116])
  );
LUT2  #(
    .INIT(4'h6)
  ) _253_ (
    .I0(ko[117]),
    .I1(ki[85]),
    .O(ko[85])
  );
LUT2  #(
    .INIT(4'h6)
  ) _254_ (
    .I0(ki[117]),
    .I1(so[21]),
    .O(ko[117])
  );
LUT2  #(
    .INIT(4'h6)
  ) _255_ (
    .I0(ko[118]),
    .I1(ki[86]),
    .O(ko[86])
  );
LUT2  #(
    .INIT(4'h6)
  ) _256_ (
    .I0(ki[118]),
    .I1(so[22]),
    .O(ko[118])
  );
LUT2  #(
    .INIT(4'h6)
  ) _257_ (
    .I0(ko[119]),
    .I1(ki[87]),
    .O(ko[87])
  );
LUT2  #(
    .INIT(4'h6)
  ) _258_ (
    .I0(ki[119]),
    .I1(so[23]),
    .O(ko[119])
  );
LUT6  #(
    .INIT(64'h07f8f807f80707f8)
  ) _259_ (
    .I0(_000_[0]),
    .I1(Rrg[8]),
    .I2(Rrg[0]),
    .I3(ki[88]),
    .I4(ki[120]),
    .I5(so[24]),
    .O(ko[88])
  );
LUT6  #(
    .INIT(64'hf10e0ef10ef1f10e)
  ) _260_ (
    .I0(_010_[0]),
    .I1(Rrg[1]),
    .I2(Rrg[0]),
    .I3(ki[89]),
    .I4(ki[121]),
    .I5(so[25]),
    .O(ko[89])
  );
LUT5  #(
    .INIT(32'd3024833460)
  ) _261_ (
    .I0(_020_[0]),
    .I1(_020_[1]),
    .I2(ki[90]),
    .I3(ki[122]),
    .I4(so[26]),
    .O(ko[90])
  );
LUT5  #(
    .INIT(32'd3024833460)
  ) _262_ (
    .I0(_023_[0]),
    .I1(_023_[1]),
    .I2(ki[91]),
    .I3(ki[123]),
    .I4(so[27]),
    .O(ko[91])
  );
LUT6  #(
    .INIT(64'h1fe0e01fe01f1fe0)
  ) _263_ (
    .I0(_026_[0]),
    .I1(Rrg[4]),
    .I2(_026_[2]),
    .I3(ki[92]),
    .I4(ki[124]),
    .I5(so[28]),
    .O(ko[92])
  );
LUT5  #(
    .INIT(32'd3024833460)
  ) _264_ (
    .I0(_035_[0]),
    .I1(_035_[1]),
    .I2(ki[93]),
    .I3(ki[125]),
    .I4(so[29]),
    .O(ko[93])
  );
LUT5  #(
    .INIT(32'd2022147960)
  ) _265_ (
    .I0(_035_[1]),
    .I1(_038_[1]),
    .I2(ki[94]),
    .I3(ki[126]),
    .I4(so[30]),
    .O(ko[94])
  );
LUT5  #(
    .INIT(32'd2022147960)
  ) _266_ (
    .I0(_035_[1]),
    .I1(_041_[1]),
    .I2(ki[95]),
    .I3(ki[127]),
    .I4(so[31]),
    .O(ko[95])
  );
LUT5  #(
    .INIT(32'd4161210360)
  ) _267_ (
    .I0(_000_[0]),
    .I1(Rrg[8]),
    .I2(Rrg[0]),
    .I3(ki[120]),
    .I4(so[24]),
    .O(ko[120])
  );
LUT5  #(
    .INIT(32'd250736910)
  ) _268_ (
    .I0(_010_[0]),
    .I1(Rrg[1]),
    .I2(Rrg[0]),
    .I3(ki[121]),
    .I4(so[25]),
    .O(ko[121])
  );
LUT4  #(
    .INIT(16'h4bb4)
  ) _269_ (
    .I0(_020_[0]),
    .I1(_020_[1]),
    .I2(ki[122]),
    .I3(so[26]),
    .O(ko[122])
  );
LUT4  #(
    .INIT(16'h4bb4)
  ) _270_ (
    .I0(_023_[0]),
    .I1(_023_[1]),
    .I2(ki[123]),
    .I3(so[27]),
    .O(ko[123])
  );
LUT5  #(
    .INIT(32'd3760136160)
  ) _271_ (
    .I0(_026_[0]),
    .I1(Rrg[4]),
    .I2(_026_[2]),
    .I3(ki[124]),
    .I4(so[28]),
    .O(ko[124])
  );
LUT4  #(
    .INIT(16'h4bb4)
  ) _272_ (
    .I0(_035_[0]),
    .I1(_035_[1]),
    .I2(ki[125]),
    .I3(so[29]),
    .O(ko[125])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _273_ (
    .I0(_035_[1]),
    .I1(_038_[1]),
    .I2(ki[126]),
    .I3(so[30]),
    .O(ko[126])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _274_ (
    .I0(_035_[1]),
    .I1(_041_[1]),
    .I2(ki[127]),
    .I3(so[31]),
    .O(ko[127])
  );
LUT4  #(
    .INIT(16'h3c5a)
  ) _275_ (
    .I0(mx[0]),
    .I1(sb[32]),
    .I2(ki[0]),
    .I3(Rrg[0]),
    .O(\do [0])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _276_ (
    .I0(sb[33]),
    .I1(mx[1]),
    .I2(Rrg[0]),
    .I3(ki[1]),
    .O(\do [1])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _277_ (
    .I0(sb[34]),
    .I1(mx[2]),
    .I2(Rrg[0]),
    .I3(ki[2]),
    .O(\do [2])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _278_ (
    .I0(sb[35]),
    .I1(mx[3]),
    .I2(Rrg[0]),
    .I3(ki[3]),
    .O(\do [3])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _279_ (
    .I0(sb[36]),
    .I1(mx[4]),
    .I2(Rrg[0]),
    .I3(ki[4]),
    .O(\do [4])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _280_ (
    .I0(sb[37]),
    .I1(mx[5]),
    .I2(Rrg[0]),
    .I3(ki[5]),
    .O(\do [5])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _281_ (
    .I0(sb[38]),
    .I1(mx[6]),
    .I2(Rrg[0]),
    .I3(ki[6]),
    .O(\do [6])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _282_ (
    .I0(sb[39]),
    .I1(mx[7]),
    .I2(Rrg[0]),
    .I3(ki[7]),
    .O(\do [7])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _283_ (
    .I0(sb[72]),
    .I1(mx[8]),
    .I2(Rrg[0]),
    .I3(ki[8]),
    .O(\do [8])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _284_ (
    .I0(sb[73]),
    .I1(mx[9]),
    .I2(Rrg[0]),
    .I3(ki[9]),
    .O(\do [9])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _285_ (
    .I0(sb[74]),
    .I1(mx[10]),
    .I2(Rrg[0]),
    .I3(ki[10]),
    .O(\do [10])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _286_ (
    .I0(sb[75]),
    .I1(mx[11]),
    .I2(Rrg[0]),
    .I3(ki[11]),
    .O(\do [11])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _287_ (
    .I0(sb[76]),
    .I1(mx[12]),
    .I2(Rrg[0]),
    .I3(ki[12]),
    .O(\do [12])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _288_ (
    .I0(sb[77]),
    .I1(mx[13]),
    .I2(Rrg[0]),
    .I3(ki[13]),
    .O(\do [13])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _289_ (
    .I0(sb[78]),
    .I1(mx[14]),
    .I2(Rrg[0]),
    .I3(ki[14]),
    .O(\do [14])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _290_ (
    .I0(sb[79]),
    .I1(mx[15]),
    .I2(Rrg[0]),
    .I3(ki[15]),
    .O(\do [15])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _291_ (
    .I0(sb[112]),
    .I1(mx[16]),
    .I2(Rrg[0]),
    .I3(ki[16]),
    .O(\do [16])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _292_ (
    .I0(sb[113]),
    .I1(mx[17]),
    .I2(Rrg[0]),
    .I3(ki[17]),
    .O(\do [17])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _293_ (
    .I0(sb[114]),
    .I1(mx[18]),
    .I2(Rrg[0]),
    .I3(ki[18]),
    .O(\do [18])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _294_ (
    .I0(sb[115]),
    .I1(mx[19]),
    .I2(Rrg[0]),
    .I3(ki[19]),
    .O(\do [19])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _295_ (
    .I0(sb[116]),
    .I1(mx[20]),
    .I2(Rrg[0]),
    .I3(ki[20]),
    .O(\do [20])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _296_ (
    .I0(sb[117]),
    .I1(mx[21]),
    .I2(Rrg[0]),
    .I3(ki[21]),
    .O(\do [21])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _297_ (
    .I0(sb[118]),
    .I1(mx[22]),
    .I2(Rrg[0]),
    .I3(ki[22]),
    .O(\do [22])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _298_ (
    .I0(sb[119]),
    .I1(mx[23]),
    .I2(Rrg[0]),
    .I3(ki[23]),
    .O(\do [23])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _299_ (
    .I0(sb[24]),
    .I1(mx[24]),
    .I2(Rrg[0]),
    .I3(ki[24]),
    .O(\do [24])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _300_ (
    .I0(sb[25]),
    .I1(mx[25]),
    .I2(Rrg[0]),
    .I3(ki[25]),
    .O(\do [25])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _301_ (
    .I0(sb[26]),
    .I1(mx[26]),
    .I2(Rrg[0]),
    .I3(ki[26]),
    .O(\do [26])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _302_ (
    .I0(sb[27]),
    .I1(mx[27]),
    .I2(Rrg[0]),
    .I3(ki[27]),
    .O(\do [27])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _303_ (
    .I0(sb[28]),
    .I1(mx[28]),
    .I2(Rrg[0]),
    .I3(ki[28]),
    .O(\do [28])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _304_ (
    .I0(sb[29]),
    .I1(mx[29]),
    .I2(Rrg[0]),
    .I3(ki[29]),
    .O(\do [29])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _305_ (
    .I0(sb[30]),
    .I1(mx[30]),
    .I2(Rrg[0]),
    .I3(ki[30]),
    .O(\do [30])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _306_ (
    .I0(sb[31]),
    .I1(mx[31]),
    .I2(Rrg[0]),
    .I3(ki[31]),
    .O(\do [31])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _307_ (
    .I0(sb[64]),
    .I1(mx[32]),
    .I2(Rrg[0]),
    .I3(ki[32]),
    .O(\do [32])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _308_ (
    .I0(sb[65]),
    .I1(mx[33]),
    .I2(Rrg[0]),
    .I3(ki[33]),
    .O(\do [33])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _309_ (
    .I0(sb[66]),
    .I1(mx[34]),
    .I2(Rrg[0]),
    .I3(ki[34]),
    .O(\do [34])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _310_ (
    .I0(sb[67]),
    .I1(mx[35]),
    .I2(Rrg[0]),
    .I3(ki[35]),
    .O(\do [35])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _311_ (
    .I0(sb[68]),
    .I1(mx[36]),
    .I2(Rrg[0]),
    .I3(ki[36]),
    .O(\do [36])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _312_ (
    .I0(sb[69]),
    .I1(mx[37]),
    .I2(Rrg[0]),
    .I3(ki[37]),
    .O(\do [37])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _313_ (
    .I0(sb[70]),
    .I1(mx[38]),
    .I2(Rrg[0]),
    .I3(ki[38]),
    .O(\do [38])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _314_ (
    .I0(sb[71]),
    .I1(mx[39]),
    .I2(Rrg[0]),
    .I3(ki[39]),
    .O(\do [39])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _315_ (
    .I0(sb[104]),
    .I1(mx[40]),
    .I2(Rrg[0]),
    .I3(ki[40]),
    .O(\do [40])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _316_ (
    .I0(sb[105]),
    .I1(mx[41]),
    .I2(Rrg[0]),
    .I3(ki[41]),
    .O(\do [41])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _317_ (
    .I0(sb[106]),
    .I1(mx[42]),
    .I2(Rrg[0]),
    .I3(ki[42]),
    .O(\do [42])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _318_ (
    .I0(sb[107]),
    .I1(mx[43]),
    .I2(Rrg[0]),
    .I3(ki[43]),
    .O(\do [43])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _319_ (
    .I0(sb[108]),
    .I1(mx[44]),
    .I2(Rrg[0]),
    .I3(ki[44]),
    .O(\do [44])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _320_ (
    .I0(sb[109]),
    .I1(mx[45]),
    .I2(Rrg[0]),
    .I3(ki[45]),
    .O(\do [45])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _321_ (
    .I0(sb[110]),
    .I1(mx[46]),
    .I2(Rrg[0]),
    .I3(ki[46]),
    .O(\do [46])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _322_ (
    .I0(sb[111]),
    .I1(mx[47]),
    .I2(Rrg[0]),
    .I3(ki[47]),
    .O(\do [47])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _323_ (
    .I0(sb[16]),
    .I1(mx[48]),
    .I2(Rrg[0]),
    .I3(ki[48]),
    .O(\do [48])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _324_ (
    .I0(sb[17]),
    .I1(mx[49]),
    .I2(Rrg[0]),
    .I3(ki[49]),
    .O(\do [49])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _325_ (
    .I0(sb[18]),
    .I1(mx[50]),
    .I2(Rrg[0]),
    .I3(ki[50]),
    .O(\do [50])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _326_ (
    .I0(sb[19]),
    .I1(mx[51]),
    .I2(Rrg[0]),
    .I3(ki[51]),
    .O(\do [51])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _327_ (
    .I0(sb[20]),
    .I1(mx[52]),
    .I2(Rrg[0]),
    .I3(ki[52]),
    .O(\do [52])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _328_ (
    .I0(sb[21]),
    .I1(mx[53]),
    .I2(Rrg[0]),
    .I3(ki[53]),
    .O(\do [53])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _329_ (
    .I0(sb[22]),
    .I1(mx[54]),
    .I2(Rrg[0]),
    .I3(ki[54]),
    .O(\do [54])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _330_ (
    .I0(sb[23]),
    .I1(mx[55]),
    .I2(Rrg[0]),
    .I3(ki[55]),
    .O(\do [55])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _331_ (
    .I0(sb[56]),
    .I1(mx[56]),
    .I2(Rrg[0]),
    .I3(ki[56]),
    .O(\do [56])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _332_ (
    .I0(sb[57]),
    .I1(mx[57]),
    .I2(Rrg[0]),
    .I3(ki[57]),
    .O(\do [57])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _333_ (
    .I0(sb[58]),
    .I1(mx[58]),
    .I2(Rrg[0]),
    .I3(ki[58]),
    .O(\do [58])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _334_ (
    .I0(sb[59]),
    .I1(mx[59]),
    .I2(Rrg[0]),
    .I3(ki[59]),
    .O(\do [59])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _335_ (
    .I0(sb[60]),
    .I1(mx[60]),
    .I2(Rrg[0]),
    .I3(ki[60]),
    .O(\do [60])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _336_ (
    .I0(sb[61]),
    .I1(mx[61]),
    .I2(Rrg[0]),
    .I3(ki[61]),
    .O(\do [61])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _337_ (
    .I0(sb[62]),
    .I1(mx[62]),
    .I2(Rrg[0]),
    .I3(ki[62]),
    .O(\do [62])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _338_ (
    .I0(sb[63]),
    .I1(mx[63]),
    .I2(Rrg[0]),
    .I3(ki[63]),
    .O(\do [63])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _339_ (
    .I0(sb[96]),
    .I1(mx[64]),
    .I2(Rrg[0]),
    .I3(ki[64]),
    .O(\do [64])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _340_ (
    .I0(sb[97]),
    .I1(mx[65]),
    .I2(Rrg[0]),
    .I3(ki[65]),
    .O(\do [65])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _341_ (
    .I0(sb[98]),
    .I1(mx[66]),
    .I2(Rrg[0]),
    .I3(ki[66]),
    .O(\do [66])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _342_ (
    .I0(sb[99]),
    .I1(mx[67]),
    .I2(Rrg[0]),
    .I3(ki[67]),
    .O(\do [67])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _343_ (
    .I0(sb[100]),
    .I1(mx[68]),
    .I2(Rrg[0]),
    .I3(ki[68]),
    .O(\do [68])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _344_ (
    .I0(sb[101]),
    .I1(mx[69]),
    .I2(Rrg[0]),
    .I3(ki[69]),
    .O(\do [69])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _345_ (
    .I0(sb[102]),
    .I1(mx[70]),
    .I2(Rrg[0]),
    .I3(ki[70]),
    .O(\do [70])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _346_ (
    .I0(sb[103]),
    .I1(mx[71]),
    .I2(Rrg[0]),
    .I3(ki[71]),
    .O(\do [71])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _347_ (
    .I0(sb[8]),
    .I1(mx[72]),
    .I2(Rrg[0]),
    .I3(ki[72]),
    .O(\do [72])
  );
AES_Comp_MixColumns  MX0 (
    .x({ sb[31:24], sb[119:112], sb[79:72], sb[39:32] }),
    .y(mx[31:0])
  );
AES_Comp_MixColumns  MX1 (
    .x({ sb[63:56], sb[23:16], sb[111:104], sb[71:64] }),
    .y(mx[63:32])
  );
AES_Comp_MixColumns  MX2 (
    .x({ sb[95:88], sb[55:48], sb[15:8], sb[103:96] }),
    .y(mx[95:64])
  );
AES_Comp_MixColumns  MX3 (
    .x({ sb[127:120], sb[87:80], sb[47:40], sb[7:0] }),
    .y(mx[127:96])
  );
AES_Comp_SubBytesComp  SB0 (
    .x(di[31:0]),
    .y(sb[31:0])
  );
AES_Comp_SubBytesComp  SB1 (
    .x(di[63:32]),
    .y(sb[63:32])
  );
AES_Comp_SubBytesComp  SB2 (
    .x(di[95:64]),
    .y(sb[95:64])
  );
AES_Comp_SubBytesComp  SB3 (
    .x(di[127:96]),
    .y(sb[127:96])
  );
AES_Comp_SubBytesComp  SBK (
    .x({ ki[23:0], ki[31:24] }),
    .y(so)
  );
assign  _010_[6:1] = { so[25], ki[121], ki[89], ki[57], Rrg[0], Rrg[1] };
assign  _000_[6:1] = { so[24], ki[120], ki[88], ki[56], Rrg[0], Rrg[8] };
assign  _035_[6:2] = { so[29], ki[125], ki[93], ki[61], ki[29] };
assign  { _038_[6:2], _038_[0] } = { so[30], ki[126], ki[94], ki[62], ki[30], _035_[1] };
assign  _020_[6:2] = { so[26], ki[122], ki[90], ki[58], ki[26] };
assign  { _041_[6:2], _041_[0] } = { so[31], ki[127], ki[95], ki[63], ki[31], _035_[1] };
assign  _023_[6:2] = { so[27], ki[123], ki[91], ki[59], ki[27] };
assign  { _026_[6:3], _026_[1] } = { so[28], ki[124], ki[92], ki[60], Rrg[4] };
assign  \rcon$func$AES_Comp.v:349$425.x  = 10'hxxx;
assign  sr = { sb[127:120], sb[87:80], sb[47:40], sb[7:0], sb[95:88], sb[55:48], sb[15:8], sb[103:96], sb[63:56], sb[23:16], sb[111:104], sb[71:64], sb[31:24], sb[119:112], sb[79:72], sb[39:32] };
endmodule
