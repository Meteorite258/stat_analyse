module AES_Comp_DEC(Kin,  Din, Dout, Krdy, Drdy, RSTn, EN, CLK, BSY, Kvld, Dvld);
wire  [6:0] _0000_;
wire  _0001_;
wire  _0002_;
wire  [6:0] _0003_;
wire  _0004_;
wire  _0005_;
wire  _0006_;
wire  _0007_;
wire  _0008_;
wire  _0009_;
wire  _0010_;
wire  _0011_;
wire  _0012_;
wire  _0013_;
wire  _0014_;
wire  _0015_;
wire  _0016_;
wire  _0017_;
wire  _0018_;
wire  _0019_;
wire  _0020_;
wire  _0021_;
wire  _0022_;
wire  _0023_;
wire  _0024_;
wire  _0025_;
wire  _0026_;
wire  _0027_;
wire  _0028_;
wire  _0029_;
wire  _0030_;
wire  _0031_;
wire  _0032_;
wire  _0033_;
wire  _0034_;
wire  _0035_;
wire  _0036_;
wire  _0037_;
wire  _0038_;
wire  _0039_;
wire  _0040_;
wire  _0041_;
wire  _0042_;
wire  _0043_;
wire  _0044_;
wire  _0045_;
wire  _0046_;
wire  _0047_;
wire  _0048_;
wire  _0049_;
wire  _0050_;
wire  _0051_;
wire  _0052_;
wire  _0053_;
wire  _0054_;
wire  _0055_;
wire  _0056_;
wire  _0057_;
wire  _0058_;
wire  _0059_;
wire  _0060_;
wire  _0061_;
wire  _0062_;
wire  _0063_;
wire  _0064_;
wire  _0065_;
wire  _0066_;
wire  _0067_;
wire  _0068_;
wire  _0069_;
wire  _0070_;
wire  _0071_;
wire  _0072_;
wire  _0073_;
wire  _0074_;
wire  _0075_;
wire  _0076_;
wire  _0077_;
wire  _0078_;
wire  _0079_;
wire  _0080_;
wire  _0081_;
wire  _0082_;
wire  _0083_;
wire  _0084_;
wire  _0085_;
wire  _0086_;
wire  _0087_;
wire  _0088_;
wire  _0089_;
wire  _0090_;
wire  _0091_;
wire  _0092_;
wire  _0093_;
wire  _0094_;
wire  _0095_;
wire  _0096_;
wire  _0097_;
wire  _0098_;
wire  _0099_;
wire  _0100_;
wire  _0101_;
wire  _0102_;
wire  _0103_;
wire  _0104_;
wire  _0105_;
wire  _0106_;
wire  _0107_;
wire  _0108_;
wire  _0109_;
wire  _0110_;
wire  _0111_;
wire  _0112_;
wire  _0113_;
wire  _0114_;
wire  _0115_;
wire  _0116_;
wire  _0117_;
wire  _0118_;
wire  _0119_;
wire  _0120_;
wire  _0121_;
wire  _0122_;
wire  _0123_;
wire  _0124_;
wire  _0125_;
wire  _0126_;
wire  _0127_;
wire  _0128_;
wire  _0129_;
wire  _0130_;
wire  _0131_;
wire  _0132_;
wire  _0133_;
wire  _0134_;
wire  _0135_;
wire  _0136_;
wire  _0137_;
wire  _0138_;
wire  _0139_;
wire  _0140_;
wire  _0141_;
wire  _0142_;
wire  _0143_;
wire  _0144_;
wire  _0145_;
wire  _0146_;
wire  _0147_;
wire  _0148_;
wire  _0149_;
wire  _0150_;
wire  _0151_;
wire  _0152_;
wire  _0153_;
wire  _0154_;
wire  _0155_;
wire  _0156_;
wire  _0157_;
wire  _0158_;
wire  _0159_;
wire  _0160_;
wire  _0161_;
wire  _0162_;
wire  _0163_;
wire  _0164_;
wire  _0165_;
wire  _0166_;
wire  _0167_;
wire  _0168_;
wire  _0169_;
wire  _0170_;
wire  _0171_;
wire  _0172_;
wire  _0173_;
wire  _0174_;
wire  _0175_;
wire  _0176_;
wire  _0177_;
wire  _0178_;
wire  _0179_;
wire  _0180_;
wire  _0181_;
wire  _0182_;
wire  _0183_;
wire  _0184_;
wire  _0185_;
wire  _0186_;
wire  _0187_;
wire  _0188_;
wire  _0189_;
wire  _0190_;
wire  _0191_;
wire  _0192_;
wire  _0193_;
wire  _0194_;
wire  _0195_;
wire  _0196_;
wire  _0197_;
wire  _0198_;
wire  _0199_;
wire  _0200_;
wire  _0201_;
wire  _0202_;
wire  _0203_;
wire  _0204_;
wire  _0205_;
wire  _0206_;
wire  _0207_;
wire  _0208_;
wire  _0209_;
wire  _0210_;
wire  _0211_;
wire  _0212_;
wire  _0213_;
wire  _0214_;
wire  _0215_;
wire  _0216_;
wire  _0217_;
wire  _0218_;
wire  _0219_;
wire  _0220_;
wire  _0221_;
wire  _0222_;
wire  _0223_;
wire  _0224_;
wire  _0225_;
wire  _0226_;
wire  _0227_;
wire  _0228_;
wire  _0229_;
wire  _0230_;
wire  _0231_;
wire  _0232_;
wire  _0233_;
wire  _0234_;
wire  _0235_;
wire  _0236_;
wire  _0237_;
wire  _0238_;
wire  _0239_;
wire  _0240_;
wire  _0241_;
wire  _0242_;
wire  _0243_;
wire  _0244_;
wire  _0245_;
wire  _0246_;
wire  _0247_;
wire  _0248_;
wire  _0249_;
wire  _0250_;
wire  _0251_;
wire  _0252_;
wire  _0253_;
wire  _0254_;
wire  _0255_;
wire  _0256_;
wire  _0257_;
wire  _0258_;
wire  _0259_;
wire  _0260_;
wire  _0261_;
wire  _0262_;
wire  _0263_;
wire  _0264_;
wire  _0265_;
wire  _0266_;
wire  _0267_;
wire  _0268_;
wire  _0269_;
wire  _0270_;
wire  _0271_;
wire  _0272_;
wire  _0273_;
wire  _0274_;
wire  _0275_;
wire  _0276_;
wire  _0277_;
wire  _0278_;
wire  _0279_;
wire  _0280_;
wire  _0281_;
wire  _0282_;
wire  _0283_;
wire  _0284_;
wire  _0285_;
wire  _0286_;
wire  _0287_;
wire  _0288_;
wire  _0289_;
wire  _0290_;
wire  _0291_;
wire  _0292_;
wire  _0293_;
wire  _0294_;
wire  _0295_;
wire  _0296_;
wire  _0297_;
wire  _0298_;
wire  _0299_;
wire  _0300_;
wire  _0301_;
wire  _0302_;
wire  _0303_;
wire  _0304_;
wire  _0305_;
wire  _0306_;
wire  _0307_;
wire  _0308_;
wire  _0309_;
wire  _0310_;
wire  _0311_;
wire  _0312_;
wire  _0313_;
wire  _0314_;
wire  _0315_;
wire  _0316_;
wire  _0317_;
wire  _0318_;
wire  _0319_;
wire  _0320_;
wire  _0321_;
wire  _0322_;
wire  _0323_;
wire  _0324_;
wire  _0325_;
wire  _0326_;
wire  _0327_;
wire  _0328_;
wire  _0329_;
wire  _0330_;
wire  _0331_;
wire  _0332_;
wire  _0333_;
wire  _0334_;
wire  _0335_;
wire  _0336_;
wire  _0337_;
wire  _0338_;
wire  _0339_;
wire  _0340_;
wire  _0341_;
wire  _0342_;
wire  _0343_;
wire  _0344_;
wire  _0345_;
wire  _0346_;
wire  _0347_;
wire  _0348_;
wire  _0349_;
wire  _0350_;
wire  _0351_;
wire  _0352_;
wire  _0353_;
wire  _0354_;
wire  _0355_;
wire  _0356_;
wire  _0357_;
wire  _0358_;
wire  _0359_;
wire  _0360_;
wire  _0361_;
wire  _0362_;
wire  _0363_;
wire  _0364_;
wire  _0365_;
wire  _0366_;
wire  _0367_;
wire  _0368_;
wire  _0369_;
wire  _0370_;
wire  _0371_;
wire  _0372_;
wire  _0373_;
wire  _0374_;
wire  _0375_;
wire  _0376_;
wire  _0377_;
wire  _0378_;
wire  _0379_;
wire  _0380_;
wire  _0381_;
wire  _0382_;
wire  _0383_;
wire  _0384_;
wire  _0385_;
wire  _0386_;
wire  _0387_;
wire  _0388_;
wire  _0389_;
wire  _0390_;
wire  _0391_;
wire  _0392_;
wire  _0393_;
wire  _0394_;
wire  _0395_;
wire  _0396_;
wire  _0397_;
wire  _0398_;
wire  _0399_;
wire  _0400_;
wire  _0401_;
wire  _0402_;
wire  _0403_;
wire  _0404_;
wire  _0405_;
wire  _0406_;
wire  _0407_;
wire  _0408_;
wire  _0409_;
wire  _0410_;
wire  _0411_;
wire  _0412_;
wire  _0413_;
wire  _0414_;
wire  _0415_;
wire  _0416_;
wire  _0417_;
wire  _0418_;
wire  _0419_;
wire  _0420_;
wire  _0421_;
wire  _0422_;
wire  _0423_;
wire  _0424_;
wire  _0425_;
wire  _0426_;
wire  _0427_;
wire  _0428_;
wire  _0429_;
wire  _0430_;
wire  _0431_;
wire  _0432_;
wire  _0433_;
wire  _0434_;
wire  _0435_;
wire  _0436_;
wire  _0437_;
wire  _0438_;
wire  _0439_;
wire  _0440_;
wire  _0441_;
wire  _0442_;
wire  _0443_;
wire  _0444_;
wire  _0445_;
wire  _0446_;
wire  _0447_;
wire  _0448_;
wire  _0449_;
wire  _0450_;
wire  _0451_;
wire  _0452_;
wire  _0453_;
wire  _0454_;
wire  _0455_;
wire  _0456_;
wire  _0457_;
wire  _0458_;
wire  _0459_;
wire  _0460_;
wire  _0461_;
wire  _0462_;
wire  _0463_;
wire  _0464_;
wire  _0465_;
wire  _0466_;
wire  _0467_;
wire  _0468_;
wire  _0469_;
wire  _0470_;
wire  _0471_;
wire  _0472_;
wire  _0473_;
wire  _0474_;
wire  _0475_;
wire  _0476_;
wire  _0477_;
wire  _0478_;
wire  _0479_;
wire  _0480_;
wire  _0481_;
wire  _0482_;
wire  _0483_;
wire  _0484_;
wire  _0485_;
wire  _0486_;
wire  _0487_;
wire  _0488_;
wire  _0489_;
wire  _0490_;
wire  _0491_;
wire  _0492_;
wire  _0493_;
wire  _0494_;
wire  _0495_;
wire  _0496_;
wire  _0497_;
wire  _0498_;
wire  _0499_;
wire  _0500_;
wire  _0501_;
wire  _0502_;
wire  _0503_;
wire  _0504_;
wire  _0505_;
wire  _0506_;
wire  _0507_;
wire  _0508_;
wire  _0509_;
wire  _0510_;
wire  _0511_;
wire  _0512_;
wire  _0513_;
wire  _0514_;
wire  _0515_;
wire  _0516_;
wire  _0517_;
wire  _0518_;
wire  _0519_;
wire  _0520_;
wire  _0521_;
wire  _0522_;
wire  _0523_;
wire  _0524_;
wire  _0525_;
wire  _0526_;
wire  _0527_;
wire  _0528_;
wire  _0529_;
wire  _0530_;
wire  _0531_;
wire  _0532_;
wire  _0533_;
wire  _0534_;
wire  _0535_;
wire  _0536_;
wire  _0537_;
wire  _0538_;
wire  _0539_;
wire  _0540_;
wire  [5:0] _0541_;
wire  [3:0] _0542_;
wire  [4:0] _0543_;
output  BSY;
wire  BSY;
wire  BSYrg;
input  CLK;
wire  CLK;
input  [127:0] Din;
wire  [127:0] Din;
wire  [127:0] Dnext;
output  [127:0] Dout;
wire  [127:0] Dout;
input  Drdy;
wire  Drdy;
wire  [127:0] Drg;
output  Dvld;
wire  Dvld;
wire  Dvldrg;
input  EN;
wire  EN;
input  [127:0] Kin;
wire  [127:0] Kin;
wire  [127:0] Knext;
input  Krdy;
wire  Krdy;
wire  [127:0] Krg;
wire  [127:0] KrgX;
output  Kvld;
wire  Kvld;
wire  Kvldrg;
input  RSTn;
wire  RSTn;
wire  [9:0] Rrg;
LUT5  #(
    .INIT(32'd2147418112)
  ) _0544_ (
    .I0(_0543_[0]),
    .I1(_0000_[2]),
    .I2(_0000_[0]),
    .I3(_0000_[1]),
    .I4(_0542_[3]),
    .O(_0008_)
  );
LUT5  #(
    .INIT(32'd4294443008)
  ) _0545_ (
    .I0(Kvldrg),
    .I1(Drdy),
    .I2(BSYrg),
    .I3(Krdy),
    .I4(EN),
    .O(_0542_[3])
  );
LUT2  #(
    .INIT(4'h4)
  ) _0546_ (
    .I0(Kvldrg),
    .I1(BSYrg),
    .O(_0543_[0])
  );
LUT2  #(
    .INIT(4'h1)
  ) _0547_ (
    .I0(Rrg[5]),
    .I1(Rrg[6]),
    .O(_0000_[2])
  );
LUT2  #(
    .INIT(4'h1)
  ) _0548_ (
    .I0(Rrg[7]),
    .I1(Rrg[8]),
    .O(_0000_[0])
  );
LUT6  #(
    .INIT(64'h0000000000000001)
  ) _0549_ (
    .I0(Rrg[9]),
    .I1(Rrg[0]),
    .I2(Rrg[1]),
    .I3(Rrg[2]),
    .I4(Rrg[3]),
    .I5(Rrg[4]),
    .O(_0000_[1])
  );
LUT5  #(
    .INIT(32'd2147483648)
  ) _0550_ (
    .I0(_0543_[0]),
    .I1(_0000_[2]),
    .I2(_0000_[0]),
    .I3(_0000_[1]),
    .I4(EN),
    .O(_0009_)
  );
LUT5  #(
    .INIT(32'd2734686208)
  ) _0551_ (
    .I0(Kvldrg),
    .I1(Krdy),
    .I2(BSYrg),
    .I3(RSTn),
    .I4(_0542_[3]),
    .O(_0010_)
  );
LUT3  #(
    .INIT(8'hd0)
  ) _0552_ (
    .I0(BSYrg),
    .I1(_0541_[2]),
    .I2(_0542_[3]),
    .O(_0006_)
  );
LUT2  #(
    .INIT(4'h8)
  ) _0553_ (
    .I0(Rrg[9]),
    .I1(Kvldrg),
    .O(_0541_[2])
  );
LUT3  #(
    .INIT(8'he0)
  ) _0554_ (
    .I0(BSYrg),
    .I1(Krdy),
    .I2(EN),
    .O(_0007_)
  );
LUT2  #(
    .INIT(4'h8)
  ) _0555_ (
    .I0(_0542_[3]),
    .I1(RSTn),
    .O(_0011_)
  );
LUT4  #(
    .INIT(16'h7000)
  ) _0556_ (
    .I0(BSYrg),
    .I1(_0541_[2]),
    .I2(RSTn),
    .I3(_0542_[3]),
    .O(_0012_)
  );
LUT1  #(
    .INIT(2'h1)
  ) _0557_ (
    .I0(_0000_[4]),
    .O(_0001_)
  );
LUT6  #(
    .INIT(64'h000000ff00007f7f)
  ) _0558_ (
    .I0(_0000_[0]),
    .I1(_0000_[1]),
    .I2(_0000_[2]),
    .I3(Rrg[9]),
    .I4(_0000_[4]),
    .I5(Kvldrg),
    .O(_0002_)
  );
MUXF7  _0559_ (
    .I0(_0001_),
    .I1(_0002_),
    .O(_0273_),
    .S(BSYrg)
  );
LUT4  #(
    .INIT(16'h0007)
  ) _0560_ (
    .I0(Drdy),
    .I1(Kvldrg),
    .I2(BSYrg),
    .I3(Krdy),
    .O(_0000_[4])
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0561_ (
    .I0(Kin[0]),
    .I1(Krg[0]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[0]),
    .I5(BSYrg),
    .O(_0275_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0562_ (
    .I0(Kin[1]),
    .I1(Krg[1]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[1]),
    .I5(BSYrg),
    .O(_0314_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0563_ (
    .I0(Kin[2]),
    .I1(Krg[2]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[2]),
    .I5(BSYrg),
    .O(_0325_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0564_ (
    .I0(Kin[3]),
    .I1(Krg[3]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[3]),
    .I5(BSYrg),
    .O(_0336_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0565_ (
    .I0(Kin[4]),
    .I1(Krg[4]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[4]),
    .I5(BSYrg),
    .O(_0347_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0566_ (
    .I0(Kin[5]),
    .I1(Krg[5]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[5]),
    .I5(BSYrg),
    .O(_0358_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0567_ (
    .I0(Kin[6]),
    .I1(Krg[6]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[6]),
    .I5(BSYrg),
    .O(_0369_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0568_ (
    .I0(Kin[7]),
    .I1(Krg[7]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[7]),
    .I5(BSYrg),
    .O(_0380_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0569_ (
    .I0(Kin[8]),
    .I1(Krg[8]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[8]),
    .I5(BSYrg),
    .O(_0391_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0570_ (
    .I0(Kin[9]),
    .I1(Krg[9]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[9]),
    .I5(BSYrg),
    .O(_0402_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0571_ (
    .I0(Kin[10]),
    .I1(Krg[10]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[10]),
    .I5(BSYrg),
    .O(_0286_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0572_ (
    .I0(Kin[11]),
    .I1(Krg[11]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[11]),
    .I5(BSYrg),
    .O(_0297_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0573_ (
    .I0(Kin[12]),
    .I1(Krg[12]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[12]),
    .I5(BSYrg),
    .O(_0306_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0574_ (
    .I0(Kin[13]),
    .I1(Krg[13]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[13]),
    .I5(BSYrg),
    .O(_0307_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0575_ (
    .I0(Kin[14]),
    .I1(Krg[14]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[14]),
    .I5(BSYrg),
    .O(_0308_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0576_ (
    .I0(Kin[15]),
    .I1(Krg[15]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[15]),
    .I5(BSYrg),
    .O(_0309_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0577_ (
    .I0(Kin[16]),
    .I1(Krg[16]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[16]),
    .I5(BSYrg),
    .O(_0310_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0578_ (
    .I0(Kin[17]),
    .I1(Krg[17]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[17]),
    .I5(BSYrg),
    .O(_0311_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0579_ (
    .I0(Kin[18]),
    .I1(Krg[18]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[18]),
    .I5(BSYrg),
    .O(_0312_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0580_ (
    .I0(Kin[19]),
    .I1(Krg[19]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[19]),
    .I5(BSYrg),
    .O(_0313_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0581_ (
    .I0(Kin[20]),
    .I1(Krg[20]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[20]),
    .I5(BSYrg),
    .O(_0315_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0582_ (
    .I0(Kin[21]),
    .I1(Krg[21]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[21]),
    .I5(BSYrg),
    .O(_0316_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0583_ (
    .I0(Kin[22]),
    .I1(Krg[22]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[22]),
    .I5(BSYrg),
    .O(_0317_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0584_ (
    .I0(Kin[23]),
    .I1(Krg[23]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[23]),
    .I5(BSYrg),
    .O(_0318_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0585_ (
    .I0(Kin[24]),
    .I1(Krg[24]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[24]),
    .I5(BSYrg),
    .O(_0319_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0586_ (
    .I0(Kin[25]),
    .I1(Krg[25]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[25]),
    .I5(BSYrg),
    .O(_0320_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0587_ (
    .I0(Kin[26]),
    .I1(Krg[26]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[26]),
    .I5(BSYrg),
    .O(_0321_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0588_ (
    .I0(Kin[27]),
    .I1(Krg[27]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[27]),
    .I5(BSYrg),
    .O(_0322_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0589_ (
    .I0(Kin[28]),
    .I1(Krg[28]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[28]),
    .I5(BSYrg),
    .O(_0323_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0590_ (
    .I0(Kin[29]),
    .I1(Krg[29]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[29]),
    .I5(BSYrg),
    .O(_0324_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0591_ (
    .I0(Kin[30]),
    .I1(Krg[30]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[30]),
    .I5(BSYrg),
    .O(_0326_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0592_ (
    .I0(Kin[31]),
    .I1(Krg[31]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[31]),
    .I5(BSYrg),
    .O(_0327_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0593_ (
    .I0(Kin[32]),
    .I1(Krg[32]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[32]),
    .I5(BSYrg),
    .O(_0328_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0594_ (
    .I0(Kin[33]),
    .I1(Krg[33]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[33]),
    .I5(BSYrg),
    .O(_0329_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0595_ (
    .I0(Kin[34]),
    .I1(Krg[34]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[34]),
    .I5(BSYrg),
    .O(_0330_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0596_ (
    .I0(Kin[35]),
    .I1(Krg[35]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[35]),
    .I5(BSYrg),
    .O(_0331_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0597_ (
    .I0(Kin[36]),
    .I1(Krg[36]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[36]),
    .I5(BSYrg),
    .O(_0332_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0598_ (
    .I0(Kin[37]),
    .I1(Krg[37]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[37]),
    .I5(BSYrg),
    .O(_0333_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0599_ (
    .I0(Kin[38]),
    .I1(Krg[38]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[38]),
    .I5(BSYrg),
    .O(_0334_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0600_ (
    .I0(Kin[39]),
    .I1(Krg[39]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[39]),
    .I5(BSYrg),
    .O(_0335_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0601_ (
    .I0(Kin[40]),
    .I1(Krg[40]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[40]),
    .I5(BSYrg),
    .O(_0337_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0602_ (
    .I0(Kin[41]),
    .I1(Krg[41]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[41]),
    .I5(BSYrg),
    .O(_0338_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0603_ (
    .I0(Kin[42]),
    .I1(Krg[42]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[42]),
    .I5(BSYrg),
    .O(_0339_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0604_ (
    .I0(Kin[43]),
    .I1(Krg[43]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[43]),
    .I5(BSYrg),
    .O(_0340_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0605_ (
    .I0(Kin[44]),
    .I1(Krg[44]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[44]),
    .I5(BSYrg),
    .O(_0341_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0606_ (
    .I0(Kin[45]),
    .I1(Krg[45]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[45]),
    .I5(BSYrg),
    .O(_0342_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0607_ (
    .I0(Kin[46]),
    .I1(Krg[46]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[46]),
    .I5(BSYrg),
    .O(_0343_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0608_ (
    .I0(Kin[47]),
    .I1(Krg[47]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[47]),
    .I5(BSYrg),
    .O(_0344_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0609_ (
    .I0(Kin[48]),
    .I1(Krg[48]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[48]),
    .I5(BSYrg),
    .O(_0345_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0610_ (
    .I0(Kin[49]),
    .I1(Krg[49]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[49]),
    .I5(BSYrg),
    .O(_0346_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0611_ (
    .I0(Kin[50]),
    .I1(Krg[50]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[50]),
    .I5(BSYrg),
    .O(_0348_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0612_ (
    .I0(Kin[51]),
    .I1(Krg[51]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[51]),
    .I5(BSYrg),
    .O(_0349_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0613_ (
    .I0(Kin[52]),
    .I1(Krg[52]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[52]),
    .I5(BSYrg),
    .O(_0350_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0614_ (
    .I0(Kin[53]),
    .I1(Krg[53]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[53]),
    .I5(BSYrg),
    .O(_0351_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0615_ (
    .I0(Kin[54]),
    .I1(Krg[54]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[54]),
    .I5(BSYrg),
    .O(_0352_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0616_ (
    .I0(Kin[55]),
    .I1(Krg[55]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[55]),
    .I5(BSYrg),
    .O(_0353_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0617_ (
    .I0(Kin[56]),
    .I1(Krg[56]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[56]),
    .I5(BSYrg),
    .O(_0354_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0618_ (
    .I0(Kin[57]),
    .I1(Krg[57]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[57]),
    .I5(BSYrg),
    .O(_0355_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0619_ (
    .I0(Kin[58]),
    .I1(Krg[58]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[58]),
    .I5(BSYrg),
    .O(_0356_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0620_ (
    .I0(Kin[59]),
    .I1(Krg[59]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[59]),
    .I5(BSYrg),
    .O(_0357_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0621_ (
    .I0(Kin[60]),
    .I1(Krg[60]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[60]),
    .I5(BSYrg),
    .O(_0359_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0622_ (
    .I0(Kin[61]),
    .I1(Krg[61]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[61]),
    .I5(BSYrg),
    .O(_0360_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0623_ (
    .I0(Kin[62]),
    .I1(Krg[62]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[62]),
    .I5(BSYrg),
    .O(_0361_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0624_ (
    .I0(Kin[63]),
    .I1(Krg[63]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[63]),
    .I5(BSYrg),
    .O(_0362_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0625_ (
    .I0(Kin[64]),
    .I1(Krg[64]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[64]),
    .I5(BSYrg),
    .O(_0363_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0626_ (
    .I0(Kin[65]),
    .I1(Krg[65]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[65]),
    .I5(BSYrg),
    .O(_0364_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0627_ (
    .I0(Kin[66]),
    .I1(Krg[66]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[66]),
    .I5(BSYrg),
    .O(_0365_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0628_ (
    .I0(Kin[67]),
    .I1(Krg[67]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[67]),
    .I5(BSYrg),
    .O(_0366_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0629_ (
    .I0(Kin[68]),
    .I1(Krg[68]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[68]),
    .I5(BSYrg),
    .O(_0367_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0630_ (
    .I0(Kin[69]),
    .I1(Krg[69]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[69]),
    .I5(BSYrg),
    .O(_0368_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0631_ (
    .I0(Kin[70]),
    .I1(Krg[70]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[70]),
    .I5(BSYrg),
    .O(_0370_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0632_ (
    .I0(Kin[71]),
    .I1(Krg[71]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[71]),
    .I5(BSYrg),
    .O(_0371_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0633_ (
    .I0(Kin[72]),
    .I1(Krg[72]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[72]),
    .I5(BSYrg),
    .O(_0372_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0634_ (
    .I0(Kin[73]),
    .I1(Krg[73]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[73]),
    .I5(BSYrg),
    .O(_0373_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0635_ (
    .I0(Kin[74]),
    .I1(Krg[74]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[74]),
    .I5(BSYrg),
    .O(_0374_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0636_ (
    .I0(Kin[75]),
    .I1(Krg[75]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[75]),
    .I5(BSYrg),
    .O(_0375_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0637_ (
    .I0(Kin[76]),
    .I1(Krg[76]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[76]),
    .I5(BSYrg),
    .O(_0376_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0638_ (
    .I0(Kin[77]),
    .I1(Krg[77]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[77]),
    .I5(BSYrg),
    .O(_0377_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0639_ (
    .I0(Kin[78]),
    .I1(Krg[78]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[78]),
    .I5(BSYrg),
    .O(_0378_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0640_ (
    .I0(Kin[79]),
    .I1(Krg[79]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[79]),
    .I5(BSYrg),
    .O(_0379_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0641_ (
    .I0(Kin[80]),
    .I1(Krg[80]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[80]),
    .I5(BSYrg),
    .O(_0381_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0642_ (
    .I0(Kin[81]),
    .I1(Krg[81]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[81]),
    .I5(BSYrg),
    .O(_0382_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0643_ (
    .I0(Kin[82]),
    .I1(Krg[82]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[82]),
    .I5(BSYrg),
    .O(_0383_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0644_ (
    .I0(Kin[83]),
    .I1(Krg[83]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[83]),
    .I5(BSYrg),
    .O(_0384_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0645_ (
    .I0(Kin[84]),
    .I1(Krg[84]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[84]),
    .I5(BSYrg),
    .O(_0385_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0646_ (
    .I0(Kin[85]),
    .I1(Krg[85]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[85]),
    .I5(BSYrg),
    .O(_0386_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0647_ (
    .I0(Kin[86]),
    .I1(Krg[86]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[86]),
    .I5(BSYrg),
    .O(_0387_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0648_ (
    .I0(Kin[87]),
    .I1(Krg[87]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[87]),
    .I5(BSYrg),
    .O(_0388_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0649_ (
    .I0(Kin[88]),
    .I1(Krg[88]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[88]),
    .I5(BSYrg),
    .O(_0389_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0650_ (
    .I0(Kin[89]),
    .I1(Krg[89]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[89]),
    .I5(BSYrg),
    .O(_0390_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0651_ (
    .I0(Kin[90]),
    .I1(Krg[90]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[90]),
    .I5(BSYrg),
    .O(_0392_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0652_ (
    .I0(Kin[91]),
    .I1(Krg[91]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[91]),
    .I5(BSYrg),
    .O(_0393_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0653_ (
    .I0(Kin[92]),
    .I1(Krg[92]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[92]),
    .I5(BSYrg),
    .O(_0394_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0654_ (
    .I0(Kin[93]),
    .I1(Krg[93]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[93]),
    .I5(BSYrg),
    .O(_0395_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0655_ (
    .I0(Kin[94]),
    .I1(Krg[94]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[94]),
    .I5(BSYrg),
    .O(_0396_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0656_ (
    .I0(Kin[95]),
    .I1(Krg[95]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[95]),
    .I5(BSYrg),
    .O(_0397_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0657_ (
    .I0(Kin[96]),
    .I1(Krg[96]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[96]),
    .I5(BSYrg),
    .O(_0398_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0658_ (
    .I0(Kin[97]),
    .I1(Krg[97]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[97]),
    .I5(BSYrg),
    .O(_0399_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0659_ (
    .I0(Kin[98]),
    .I1(Krg[98]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[98]),
    .I5(BSYrg),
    .O(_0400_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0660_ (
    .I0(Kin[99]),
    .I1(Krg[99]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[99]),
    .I5(BSYrg),
    .O(_0401_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0661_ (
    .I0(Kin[100]),
    .I1(Krg[100]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[100]),
    .I5(BSYrg),
    .O(_0276_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0662_ (
    .I0(Kin[101]),
    .I1(Krg[101]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[101]),
    .I5(BSYrg),
    .O(_0277_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0663_ (
    .I0(Kin[102]),
    .I1(Krg[102]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[102]),
    .I5(BSYrg),
    .O(_0278_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0664_ (
    .I0(Kin[103]),
    .I1(Krg[103]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[103]),
    .I5(BSYrg),
    .O(_0279_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0665_ (
    .I0(Kin[104]),
    .I1(Krg[104]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[104]),
    .I5(BSYrg),
    .O(_0280_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0666_ (
    .I0(Kin[105]),
    .I1(Krg[105]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[105]),
    .I5(BSYrg),
    .O(_0281_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0667_ (
    .I0(Kin[106]),
    .I1(Krg[106]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[106]),
    .I5(BSYrg),
    .O(_0282_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0668_ (
    .I0(Kin[107]),
    .I1(Krg[107]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[107]),
    .I5(BSYrg),
    .O(_0283_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0669_ (
    .I0(Kin[108]),
    .I1(Krg[108]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[108]),
    .I5(BSYrg),
    .O(_0284_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0670_ (
    .I0(Kin[109]),
    .I1(Krg[109]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[109]),
    .I5(BSYrg),
    .O(_0285_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0671_ (
    .I0(Kin[110]),
    .I1(Krg[110]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[110]),
    .I5(BSYrg),
    .O(_0287_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0672_ (
    .I0(Kin[111]),
    .I1(Krg[111]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[111]),
    .I5(BSYrg),
    .O(_0288_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0673_ (
    .I0(Kin[112]),
    .I1(Krg[112]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[112]),
    .I5(BSYrg),
    .O(_0289_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0674_ (
    .I0(Kin[113]),
    .I1(Krg[113]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[113]),
    .I5(BSYrg),
    .O(_0290_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0675_ (
    .I0(Kin[114]),
    .I1(Krg[114]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[114]),
    .I5(BSYrg),
    .O(_0291_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0676_ (
    .I0(Kin[115]),
    .I1(Krg[115]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[115]),
    .I5(BSYrg),
    .O(_0292_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0677_ (
    .I0(Kin[116]),
    .I1(Krg[116]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[116]),
    .I5(BSYrg),
    .O(_0293_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0678_ (
    .I0(Kin[117]),
    .I1(Krg[117]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[117]),
    .I5(BSYrg),
    .O(_0294_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0679_ (
    .I0(Kin[118]),
    .I1(Krg[118]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[118]),
    .I5(BSYrg),
    .O(_0295_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0680_ (
    .I0(Kin[119]),
    .I1(Krg[119]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[119]),
    .I5(BSYrg),
    .O(_0296_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0681_ (
    .I0(Kin[120]),
    .I1(Krg[120]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[120]),
    .I5(BSYrg),
    .O(_0298_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0682_ (
    .I0(Kin[121]),
    .I1(Krg[121]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[121]),
    .I5(BSYrg),
    .O(_0299_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0683_ (
    .I0(Kin[122]),
    .I1(Krg[122]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[122]),
    .I5(BSYrg),
    .O(_0300_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0684_ (
    .I0(Kin[123]),
    .I1(Krg[123]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[123]),
    .I5(BSYrg),
    .O(_0301_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0685_ (
    .I0(Kin[124]),
    .I1(Krg[124]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[124]),
    .I5(BSYrg),
    .O(_0302_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0686_ (
    .I0(Kin[125]),
    .I1(Krg[125]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[125]),
    .I5(BSYrg),
    .O(_0303_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0687_ (
    .I0(Kin[126]),
    .I1(Krg[126]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[126]),
    .I5(BSYrg),
    .O(_0304_)
  );
LUT6  #(
    .INIT(64'hcfcfc0c0aaffaa00)
  ) _0688_ (
    .I0(Kin[127]),
    .I1(Krg[127]),
    .I2(_0541_[2]),
    .I3(Krdy),
    .I4(Knext[127]),
    .I5(BSYrg),
    .O(_0305_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0689_ (
    .I0(Dnext[0]),
    .I1(Krg[0]),
    .I2(Din[0]),
    .I3(BSYrg),
    .O(_0403_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0690_ (
    .I0(Dnext[1]),
    .I1(Krg[1]),
    .I2(Din[1]),
    .I3(BSYrg),
    .O(_0442_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0691_ (
    .I0(Dnext[2]),
    .I1(Krg[2]),
    .I2(Din[2]),
    .I3(BSYrg),
    .O(_0453_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0692_ (
    .I0(Dnext[3]),
    .I1(Krg[3]),
    .I2(Din[3]),
    .I3(BSYrg),
    .O(_0464_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0693_ (
    .I0(Dnext[4]),
    .I1(Krg[4]),
    .I2(Din[4]),
    .I3(BSYrg),
    .O(_0475_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0694_ (
    .I0(Dnext[5]),
    .I1(Krg[5]),
    .I2(Din[5]),
    .I3(BSYrg),
    .O(_0486_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0695_ (
    .I0(Dnext[6]),
    .I1(Krg[6]),
    .I2(Din[6]),
    .I3(BSYrg),
    .O(_0497_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0696_ (
    .I0(Dnext[7]),
    .I1(Krg[7]),
    .I2(Din[7]),
    .I3(BSYrg),
    .O(_0508_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0697_ (
    .I0(Dnext[8]),
    .I1(Krg[8]),
    .I2(Din[8]),
    .I3(BSYrg),
    .O(_0519_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0698_ (
    .I0(Dnext[9]),
    .I1(Krg[9]),
    .I2(Din[9]),
    .I3(BSYrg),
    .O(_0530_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0699_ (
    .I0(Dnext[10]),
    .I1(Krg[10]),
    .I2(Din[10]),
    .I3(BSYrg),
    .O(_0414_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0700_ (
    .I0(Dnext[11]),
    .I1(Krg[11]),
    .I2(Din[11]),
    .I3(BSYrg),
    .O(_0425_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0701_ (
    .I0(Dnext[12]),
    .I1(Krg[12]),
    .I2(Din[12]),
    .I3(BSYrg),
    .O(_0434_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0702_ (
    .I0(Dnext[13]),
    .I1(Krg[13]),
    .I2(Din[13]),
    .I3(BSYrg),
    .O(_0435_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0703_ (
    .I0(Dnext[14]),
    .I1(Krg[14]),
    .I2(Din[14]),
    .I3(BSYrg),
    .O(_0436_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0704_ (
    .I0(Dnext[15]),
    .I1(Krg[15]),
    .I2(Din[15]),
    .I3(BSYrg),
    .O(_0437_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0705_ (
    .I0(Dnext[16]),
    .I1(Krg[16]),
    .I2(Din[16]),
    .I3(BSYrg),
    .O(_0438_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0706_ (
    .I0(Dnext[17]),
    .I1(Krg[17]),
    .I2(Din[17]),
    .I3(BSYrg),
    .O(_0439_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0707_ (
    .I0(Dnext[18]),
    .I1(Krg[18]),
    .I2(Din[18]),
    .I3(BSYrg),
    .O(_0440_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0708_ (
    .I0(Dnext[19]),
    .I1(Krg[19]),
    .I2(Din[19]),
    .I3(BSYrg),
    .O(_0441_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0709_ (
    .I0(Dnext[20]),
    .I1(Krg[20]),
    .I2(Din[20]),
    .I3(BSYrg),
    .O(_0443_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0710_ (
    .I0(Dnext[21]),
    .I1(Krg[21]),
    .I2(Din[21]),
    .I3(BSYrg),
    .O(_0444_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0711_ (
    .I0(Dnext[22]),
    .I1(Krg[22]),
    .I2(Din[22]),
    .I3(BSYrg),
    .O(_0445_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0712_ (
    .I0(Dnext[23]),
    .I1(Krg[23]),
    .I2(Din[23]),
    .I3(BSYrg),
    .O(_0446_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0713_ (
    .I0(Dnext[24]),
    .I1(Krg[24]),
    .I2(Din[24]),
    .I3(BSYrg),
    .O(_0447_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0714_ (
    .I0(Dnext[25]),
    .I1(Krg[25]),
    .I2(Din[25]),
    .I3(BSYrg),
    .O(_0448_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0715_ (
    .I0(Dnext[26]),
    .I1(Krg[26]),
    .I2(Din[26]),
    .I3(BSYrg),
    .O(_0449_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0716_ (
    .I0(Dnext[27]),
    .I1(Krg[27]),
    .I2(Din[27]),
    .I3(BSYrg),
    .O(_0450_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0717_ (
    .I0(Dnext[28]),
    .I1(Krg[28]),
    .I2(Din[28]),
    .I3(BSYrg),
    .O(_0451_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0718_ (
    .I0(Dnext[29]),
    .I1(Krg[29]),
    .I2(Din[29]),
    .I3(BSYrg),
    .O(_0452_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0719_ (
    .I0(Dnext[30]),
    .I1(Krg[30]),
    .I2(Din[30]),
    .I3(BSYrg),
    .O(_0454_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0720_ (
    .I0(Dnext[31]),
    .I1(Krg[31]),
    .I2(Din[31]),
    .I3(BSYrg),
    .O(_0455_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0721_ (
    .I0(Dnext[32]),
    .I1(Krg[32]),
    .I2(Din[32]),
    .I3(BSYrg),
    .O(_0456_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0722_ (
    .I0(Dnext[33]),
    .I1(Krg[33]),
    .I2(Din[33]),
    .I3(BSYrg),
    .O(_0457_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0723_ (
    .I0(Dnext[34]),
    .I1(Krg[34]),
    .I2(Din[34]),
    .I3(BSYrg),
    .O(_0458_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0724_ (
    .I0(Dnext[35]),
    .I1(Krg[35]),
    .I2(Din[35]),
    .I3(BSYrg),
    .O(_0459_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0725_ (
    .I0(Dnext[36]),
    .I1(Krg[36]),
    .I2(Din[36]),
    .I3(BSYrg),
    .O(_0460_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0726_ (
    .I0(Dnext[37]),
    .I1(Krg[37]),
    .I2(Din[37]),
    .I3(BSYrg),
    .O(_0461_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0727_ (
    .I0(Dnext[38]),
    .I1(Krg[38]),
    .I2(Din[38]),
    .I3(BSYrg),
    .O(_0462_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0728_ (
    .I0(Dnext[39]),
    .I1(Krg[39]),
    .I2(Din[39]),
    .I3(BSYrg),
    .O(_0463_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0729_ (
    .I0(Dnext[40]),
    .I1(Krg[40]),
    .I2(Din[40]),
    .I3(BSYrg),
    .O(_0465_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0730_ (
    .I0(Dnext[41]),
    .I1(Krg[41]),
    .I2(Din[41]),
    .I3(BSYrg),
    .O(_0466_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0731_ (
    .I0(Dnext[42]),
    .I1(Krg[42]),
    .I2(Din[42]),
    .I3(BSYrg),
    .O(_0467_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0732_ (
    .I0(Dnext[43]),
    .I1(Krg[43]),
    .I2(Din[43]),
    .I3(BSYrg),
    .O(_0468_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0733_ (
    .I0(Dnext[44]),
    .I1(Krg[44]),
    .I2(Din[44]),
    .I3(BSYrg),
    .O(_0469_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0734_ (
    .I0(Dnext[45]),
    .I1(Krg[45]),
    .I2(Din[45]),
    .I3(BSYrg),
    .O(_0470_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0735_ (
    .I0(Dnext[46]),
    .I1(Krg[46]),
    .I2(Din[46]),
    .I3(BSYrg),
    .O(_0471_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0736_ (
    .I0(Dnext[47]),
    .I1(Krg[47]),
    .I2(Din[47]),
    .I3(BSYrg),
    .O(_0472_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0737_ (
    .I0(Dnext[48]),
    .I1(Krg[48]),
    .I2(Din[48]),
    .I3(BSYrg),
    .O(_0473_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0738_ (
    .I0(Dnext[49]),
    .I1(Krg[49]),
    .I2(Din[49]),
    .I3(BSYrg),
    .O(_0474_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0739_ (
    .I0(Dnext[50]),
    .I1(Krg[50]),
    .I2(Din[50]),
    .I3(BSYrg),
    .O(_0476_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0740_ (
    .I0(Dnext[51]),
    .I1(Krg[51]),
    .I2(Din[51]),
    .I3(BSYrg),
    .O(_0477_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0741_ (
    .I0(Dnext[52]),
    .I1(Krg[52]),
    .I2(Din[52]),
    .I3(BSYrg),
    .O(_0478_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0742_ (
    .I0(Dnext[53]),
    .I1(Krg[53]),
    .I2(Din[53]),
    .I3(BSYrg),
    .O(_0479_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0743_ (
    .I0(Dnext[54]),
    .I1(Krg[54]),
    .I2(Din[54]),
    .I3(BSYrg),
    .O(_0480_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0744_ (
    .I0(Dnext[55]),
    .I1(Krg[55]),
    .I2(Din[55]),
    .I3(BSYrg),
    .O(_0481_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0745_ (
    .I0(Dnext[56]),
    .I1(Krg[56]),
    .I2(Din[56]),
    .I3(BSYrg),
    .O(_0482_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0746_ (
    .I0(Dnext[57]),
    .I1(Krg[57]),
    .I2(Din[57]),
    .I3(BSYrg),
    .O(_0483_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0747_ (
    .I0(Dnext[58]),
    .I1(Krg[58]),
    .I2(Din[58]),
    .I3(BSYrg),
    .O(_0484_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0748_ (
    .I0(Dnext[59]),
    .I1(Krg[59]),
    .I2(Din[59]),
    .I3(BSYrg),
    .O(_0485_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0749_ (
    .I0(Dnext[60]),
    .I1(Krg[60]),
    .I2(Din[60]),
    .I3(BSYrg),
    .O(_0487_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0750_ (
    .I0(Dnext[61]),
    .I1(Krg[61]),
    .I2(Din[61]),
    .I3(BSYrg),
    .O(_0488_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0751_ (
    .I0(Dnext[62]),
    .I1(Krg[62]),
    .I2(Din[62]),
    .I3(BSYrg),
    .O(_0489_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0752_ (
    .I0(Dnext[63]),
    .I1(Krg[63]),
    .I2(Din[63]),
    .I3(BSYrg),
    .O(_0490_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0753_ (
    .I0(Dnext[64]),
    .I1(Krg[64]),
    .I2(Din[64]),
    .I3(BSYrg),
    .O(_0491_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0754_ (
    .I0(Dnext[65]),
    .I1(Krg[65]),
    .I2(Din[65]),
    .I3(BSYrg),
    .O(_0492_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0755_ (
    .I0(Dnext[66]),
    .I1(Krg[66]),
    .I2(Din[66]),
    .I3(BSYrg),
    .O(_0493_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0756_ (
    .I0(Dnext[67]),
    .I1(Krg[67]),
    .I2(Din[67]),
    .I3(BSYrg),
    .O(_0494_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0757_ (
    .I0(Dnext[68]),
    .I1(Krg[68]),
    .I2(Din[68]),
    .I3(BSYrg),
    .O(_0495_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0758_ (
    .I0(Dnext[69]),
    .I1(Krg[69]),
    .I2(Din[69]),
    .I3(BSYrg),
    .O(_0496_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0759_ (
    .I0(Dnext[70]),
    .I1(Krg[70]),
    .I2(Din[70]),
    .I3(BSYrg),
    .O(_0498_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0760_ (
    .I0(Dnext[71]),
    .I1(Krg[71]),
    .I2(Din[71]),
    .I3(BSYrg),
    .O(_0499_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0761_ (
    .I0(Dnext[72]),
    .I1(Krg[72]),
    .I2(Din[72]),
    .I3(BSYrg),
    .O(_0500_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0762_ (
    .I0(Dnext[73]),
    .I1(Krg[73]),
    .I2(Din[73]),
    .I3(BSYrg),
    .O(_0501_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0763_ (
    .I0(Dnext[74]),
    .I1(Krg[74]),
    .I2(Din[74]),
    .I3(BSYrg),
    .O(_0502_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0764_ (
    .I0(Dnext[75]),
    .I1(Krg[75]),
    .I2(Din[75]),
    .I3(BSYrg),
    .O(_0503_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0765_ (
    .I0(Dnext[76]),
    .I1(Krg[76]),
    .I2(Din[76]),
    .I3(BSYrg),
    .O(_0504_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0766_ (
    .I0(Dnext[77]),
    .I1(Krg[77]),
    .I2(Din[77]),
    .I3(BSYrg),
    .O(_0505_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0767_ (
    .I0(Dnext[78]),
    .I1(Krg[78]),
    .I2(Din[78]),
    .I3(BSYrg),
    .O(_0506_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0768_ (
    .I0(Dnext[79]),
    .I1(Krg[79]),
    .I2(Din[79]),
    .I3(BSYrg),
    .O(_0507_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0769_ (
    .I0(Dnext[80]),
    .I1(Krg[80]),
    .I2(Din[80]),
    .I3(BSYrg),
    .O(_0509_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0770_ (
    .I0(Dnext[81]),
    .I1(Krg[81]),
    .I2(Din[81]),
    .I3(BSYrg),
    .O(_0510_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0771_ (
    .I0(Dnext[82]),
    .I1(Krg[82]),
    .I2(Din[82]),
    .I3(BSYrg),
    .O(_0511_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0772_ (
    .I0(Dnext[83]),
    .I1(Krg[83]),
    .I2(Din[83]),
    .I3(BSYrg),
    .O(_0512_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0773_ (
    .I0(Dnext[84]),
    .I1(Krg[84]),
    .I2(Din[84]),
    .I3(BSYrg),
    .O(_0513_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0774_ (
    .I0(Dnext[85]),
    .I1(Krg[85]),
    .I2(Din[85]),
    .I3(BSYrg),
    .O(_0514_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0775_ (
    .I0(Dnext[86]),
    .I1(Krg[86]),
    .I2(Din[86]),
    .I3(BSYrg),
    .O(_0515_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0776_ (
    .I0(Dnext[87]),
    .I1(Krg[87]),
    .I2(Din[87]),
    .I3(BSYrg),
    .O(_0516_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0777_ (
    .I0(Dnext[88]),
    .I1(Krg[88]),
    .I2(Din[88]),
    .I3(BSYrg),
    .O(_0517_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0778_ (
    .I0(Dnext[89]),
    .I1(Krg[89]),
    .I2(Din[89]),
    .I3(BSYrg),
    .O(_0518_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0779_ (
    .I0(Dnext[90]),
    .I1(Krg[90]),
    .I2(Din[90]),
    .I3(BSYrg),
    .O(_0520_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0780_ (
    .I0(Dnext[91]),
    .I1(Krg[91]),
    .I2(Din[91]),
    .I3(BSYrg),
    .O(_0521_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0781_ (
    .I0(Dnext[92]),
    .I1(Krg[92]),
    .I2(Din[92]),
    .I3(BSYrg),
    .O(_0522_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0782_ (
    .I0(Dnext[93]),
    .I1(Krg[93]),
    .I2(Din[93]),
    .I3(BSYrg),
    .O(_0523_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0783_ (
    .I0(Dnext[94]),
    .I1(Krg[94]),
    .I2(Din[94]),
    .I3(BSYrg),
    .O(_0524_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0784_ (
    .I0(Dnext[95]),
    .I1(Krg[95]),
    .I2(Din[95]),
    .I3(BSYrg),
    .O(_0525_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0785_ (
    .I0(Dnext[96]),
    .I1(Krg[96]),
    .I2(Din[96]),
    .I3(BSYrg),
    .O(_0526_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0786_ (
    .I0(Dnext[97]),
    .I1(Krg[97]),
    .I2(Din[97]),
    .I3(BSYrg),
    .O(_0527_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0787_ (
    .I0(Dnext[98]),
    .I1(Krg[98]),
    .I2(Din[98]),
    .I3(BSYrg),
    .O(_0528_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0788_ (
    .I0(Dnext[99]),
    .I1(Krg[99]),
    .I2(Din[99]),
    .I3(BSYrg),
    .O(_0529_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0789_ (
    .I0(Dnext[100]),
    .I1(Krg[100]),
    .I2(Din[100]),
    .I3(BSYrg),
    .O(_0404_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0790_ (
    .I0(Dnext[101]),
    .I1(Krg[101]),
    .I2(Din[101]),
    .I3(BSYrg),
    .O(_0405_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0791_ (
    .I0(Dnext[102]),
    .I1(Krg[102]),
    .I2(Din[102]),
    .I3(BSYrg),
    .O(_0406_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0792_ (
    .I0(Dnext[103]),
    .I1(Krg[103]),
    .I2(Din[103]),
    .I3(BSYrg),
    .O(_0407_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0793_ (
    .I0(Dnext[104]),
    .I1(Krg[104]),
    .I2(Din[104]),
    .I3(BSYrg),
    .O(_0408_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0794_ (
    .I0(Dnext[105]),
    .I1(Krg[105]),
    .I2(Din[105]),
    .I3(BSYrg),
    .O(_0409_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0795_ (
    .I0(Dnext[106]),
    .I1(Krg[106]),
    .I2(Din[106]),
    .I3(BSYrg),
    .O(_0410_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0796_ (
    .I0(Dnext[107]),
    .I1(Krg[107]),
    .I2(Din[107]),
    .I3(BSYrg),
    .O(_0411_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0797_ (
    .I0(Dnext[108]),
    .I1(Krg[108]),
    .I2(Din[108]),
    .I3(BSYrg),
    .O(_0412_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0798_ (
    .I0(Dnext[109]),
    .I1(Krg[109]),
    .I2(Din[109]),
    .I3(BSYrg),
    .O(_0413_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0799_ (
    .I0(Dnext[110]),
    .I1(Krg[110]),
    .I2(Din[110]),
    .I3(BSYrg),
    .O(_0415_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0800_ (
    .I0(Dnext[111]),
    .I1(Krg[111]),
    .I2(Din[111]),
    .I3(BSYrg),
    .O(_0416_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0801_ (
    .I0(Dnext[112]),
    .I1(Krg[112]),
    .I2(Din[112]),
    .I3(BSYrg),
    .O(_0417_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0802_ (
    .I0(Dnext[113]),
    .I1(Krg[113]),
    .I2(Din[113]),
    .I3(BSYrg),
    .O(_0418_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0803_ (
    .I0(Dnext[114]),
    .I1(Krg[114]),
    .I2(Din[114]),
    .I3(BSYrg),
    .O(_0419_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0804_ (
    .I0(Dnext[115]),
    .I1(Krg[115]),
    .I2(Din[115]),
    .I3(BSYrg),
    .O(_0420_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0805_ (
    .I0(Dnext[116]),
    .I1(Krg[116]),
    .I2(Din[116]),
    .I3(BSYrg),
    .O(_0421_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0806_ (
    .I0(Dnext[117]),
    .I1(Krg[117]),
    .I2(Din[117]),
    .I3(BSYrg),
    .O(_0422_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0807_ (
    .I0(Dnext[118]),
    .I1(Krg[118]),
    .I2(Din[118]),
    .I3(BSYrg),
    .O(_0423_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0808_ (
    .I0(Dnext[119]),
    .I1(Krg[119]),
    .I2(Din[119]),
    .I3(BSYrg),
    .O(_0424_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0809_ (
    .I0(Dnext[120]),
    .I1(Krg[120]),
    .I2(Din[120]),
    .I3(BSYrg),
    .O(_0426_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0810_ (
    .I0(Dnext[121]),
    .I1(Krg[121]),
    .I2(Din[121]),
    .I3(BSYrg),
    .O(_0427_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0811_ (
    .I0(Dnext[122]),
    .I1(Krg[122]),
    .I2(Din[122]),
    .I3(BSYrg),
    .O(_0428_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0812_ (
    .I0(Dnext[123]),
    .I1(Krg[123]),
    .I2(Din[123]),
    .I3(BSYrg),
    .O(_0429_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0813_ (
    .I0(Dnext[124]),
    .I1(Krg[124]),
    .I2(Din[124]),
    .I3(BSYrg),
    .O(_0430_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0814_ (
    .I0(Dnext[125]),
    .I1(Krg[125]),
    .I2(Din[125]),
    .I3(BSYrg),
    .O(_0431_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0815_ (
    .I0(Dnext[126]),
    .I1(Krg[126]),
    .I2(Din[126]),
    .I3(BSYrg),
    .O(_0432_)
  );
LUT4  #(
    .INIT(16'haa3c)
  ) _0816_ (
    .I0(Dnext[127]),
    .I1(Krg[127]),
    .I2(Din[127]),
    .I3(BSYrg),
    .O(_0433_)
  );
LUT4  #(
    .INIT(16'haf0c)
  ) _0817_ (
    .I0(Kvldrg),
    .I1(Krdy),
    .I2(BSYrg),
    .I3(Rrg[1]),
    .O(_0531_)
  );
LUT5  #(
    .INIT(32'd4037685296)
  ) _0818_ (
    .I0(Rrg[0]),
    .I1(Krdy),
    .I2(Rrg[2]),
    .I3(Kvldrg),
    .I4(BSYrg),
    .O(_0532_)
  );
LUT5  #(
    .INIT(32'd4037685296)
  ) _0819_ (
    .I0(Rrg[1]),
    .I1(Krdy),
    .I2(Rrg[3]),
    .I3(Kvldrg),
    .I4(BSYrg),
    .O(_0533_)
  );
LUT5  #(
    .INIT(32'd4037685296)
  ) _0820_ (
    .I0(Rrg[2]),
    .I1(Krdy),
    .I2(Rrg[4]),
    .I3(Kvldrg),
    .I4(BSYrg),
    .O(_0534_)
  );
LUT5  #(
    .INIT(32'd4037685296)
  ) _0821_ (
    .I0(Rrg[3]),
    .I1(Krdy),
    .I2(Rrg[5]),
    .I3(Kvldrg),
    .I4(BSYrg),
    .O(_0535_)
  );
LUT5  #(
    .INIT(32'd4037685296)
  ) _0822_ (
    .I0(Rrg[4]),
    .I1(Krdy),
    .I2(Rrg[6]),
    .I3(Kvldrg),
    .I4(BSYrg),
    .O(_0536_)
  );
LUT5  #(
    .INIT(32'd4037685296)
  ) _0823_ (
    .I0(Rrg[5]),
    .I1(Krdy),
    .I2(Rrg[7]),
    .I3(Kvldrg),
    .I4(BSYrg),
    .O(_0537_)
  );
LUT5  #(
    .INIT(32'd4037685296)
  ) _0824_ (
    .I0(Rrg[6]),
    .I1(Krdy),
    .I2(Rrg[8]),
    .I3(Kvldrg),
    .I4(BSYrg),
    .O(_0538_)
  );
LUT5  #(
    .INIT(32'd1145310976)
  ) _0825_ (
    .I0(Kvldrg),
    .I1(Rrg[7]),
    .I2(Krdy),
    .I3(Rrg[9]),
    .I4(BSYrg),
    .O(_0539_)
  );
LUT1  #(
    .INIT(2'h2)
  ) _0826_ (
    .I0(_0003_[5]),
    .O(_0004_)
  );
LUT6  #(
    .INIT(64'hffffffffffffff40)
  ) _0827_ (
    .I0(Rrg[7]),
    .I1(_0000_[1]),
    .I2(_0000_[2]),
    .I3(Rrg[8]),
    .I4(Kvldrg),
    .I5(_0003_[5]),
    .O(_0005_)
  );
MUXF7  _0828_ (
    .I0(_0004_),
    .I1(_0005_),
    .O(_0540_),
    .S(_0003_[6])
  );
LUT3  #(
    .INIT(8'h10)
  ) _0829_ (
    .I0(Krdy),
    .I1(BSYrg),
    .I2(Rrg[0]),
    .O(_0003_[5])
  );
LUT4  #(
    .INIT(16'hef00)
  ) _0830_ (
    .I0(Rrg[9]),
    .I1(Rrg[0]),
    .I2(Kvldrg),
    .I3(BSYrg),
    .O(_0003_[6])
  );
LUT5  #(
    .INIT(32'd4286578688)
  ) _0831_ (
    .I0(_0000_[0]),
    .I1(_0000_[1]),
    .I2(_0000_[2]),
    .I3(Kvldrg),
    .I4(BSYrg),
    .O(_0274_)
  );
INV  _0832_ (
    .I(RSTn),
    .O(_0014_)
  );
INV  _0833_ (
    .I(Kvldrg),
    .O(_0013_)
  );
INV  _0834_ (
    .I(RSTn),
    .O(_0015_)
  );
INV  _0835_ (
    .I(RSTn),
    .O(_0016_)
  );
INV  _0836_ (
    .I(RSTn),
    .O(_0017_)
  );
INV  _0837_ (
    .I(RSTn),
    .O(_0018_)
  );
INV  _0838_ (
    .I(RSTn),
    .O(_0019_)
  );
INV  _0839_ (
    .I(RSTn),
    .O(_0020_)
  );
INV  _0840_ (
    .I(RSTn),
    .O(_0021_)
  );
INV  _0841_ (
    .I(RSTn),
    .O(_0022_)
  );
INV  _0842_ (
    .I(RSTn),
    .O(_0023_)
  );
INV  _0843_ (
    .I(RSTn),
    .O(_0024_)
  );
INV  _0844_ (
    .I(RSTn),
    .O(_0025_)
  );
INV  _0845_ (
    .I(RSTn),
    .O(_0026_)
  );
INV  _0846_ (
    .I(RSTn),
    .O(_0027_)
  );
INV  _0847_ (
    .I(RSTn),
    .O(_0028_)
  );
INV  _0848_ (
    .I(RSTn),
    .O(_0029_)
  );
INV  _0849_ (
    .I(RSTn),
    .O(_0030_)
  );
INV  _0850_ (
    .I(RSTn),
    .O(_0031_)
  );
INV  _0851_ (
    .I(RSTn),
    .O(_0032_)
  );
INV  _0852_ (
    .I(RSTn),
    .O(_0033_)
  );
INV  _0853_ (
    .I(RSTn),
    .O(_0034_)
  );
INV  _0854_ (
    .I(RSTn),
    .O(_0035_)
  );
INV  _0855_ (
    .I(RSTn),
    .O(_0036_)
  );
INV  _0856_ (
    .I(RSTn),
    .O(_0037_)
  );
INV  _0857_ (
    .I(RSTn),
    .O(_0038_)
  );
INV  _0858_ (
    .I(RSTn),
    .O(_0039_)
  );
INV  _0859_ (
    .I(RSTn),
    .O(_0040_)
  );
INV  _0860_ (
    .I(RSTn),
    .O(_0041_)
  );
INV  _0861_ (
    .I(RSTn),
    .O(_0042_)
  );
INV  _0862_ (
    .I(RSTn),
    .O(_0043_)
  );
INV  _0863_ (
    .I(RSTn),
    .O(_0044_)
  );
INV  _0864_ (
    .I(RSTn),
    .O(_0045_)
  );
INV  _0865_ (
    .I(RSTn),
    .O(_0046_)
  );
INV  _0866_ (
    .I(RSTn),
    .O(_0047_)
  );
INV  _0867_ (
    .I(RSTn),
    .O(_0048_)
  );
INV  _0868_ (
    .I(RSTn),
    .O(_0049_)
  );
INV  _0869_ (
    .I(RSTn),
    .O(_0050_)
  );
INV  _0870_ (
    .I(RSTn),
    .O(_0051_)
  );
INV  _0871_ (
    .I(RSTn),
    .O(_0052_)
  );
INV  _0872_ (
    .I(RSTn),
    .O(_0053_)
  );
INV  _0873_ (
    .I(RSTn),
    .O(_0054_)
  );
INV  _0874_ (
    .I(RSTn),
    .O(_0055_)
  );
INV  _0875_ (
    .I(RSTn),
    .O(_0056_)
  );
INV  _0876_ (
    .I(RSTn),
    .O(_0057_)
  );
INV  _0877_ (
    .I(RSTn),
    .O(_0058_)
  );
INV  _0878_ (
    .I(RSTn),
    .O(_0059_)
  );
INV  _0879_ (
    .I(RSTn),
    .O(_0060_)
  );
INV  _0880_ (
    .I(RSTn),
    .O(_0061_)
  );
INV  _0881_ (
    .I(RSTn),
    .O(_0062_)
  );
INV  _0882_ (
    .I(RSTn),
    .O(_0063_)
  );
INV  _0883_ (
    .I(RSTn),
    .O(_0064_)
  );
INV  _0884_ (
    .I(RSTn),
    .O(_0065_)
  );
INV  _0885_ (
    .I(RSTn),
    .O(_0066_)
  );
INV  _0886_ (
    .I(RSTn),
    .O(_0067_)
  );
INV  _0887_ (
    .I(RSTn),
    .O(_0068_)
  );
INV  _0888_ (
    .I(RSTn),
    .O(_0069_)
  );
INV  _0889_ (
    .I(RSTn),
    .O(_0070_)
  );
INV  _0890_ (
    .I(RSTn),
    .O(_0071_)
  );
INV  _0891_ (
    .I(RSTn),
    .O(_0072_)
  );
INV  _0892_ (
    .I(RSTn),
    .O(_0073_)
  );
INV  _0893_ (
    .I(RSTn),
    .O(_0074_)
  );
INV  _0894_ (
    .I(RSTn),
    .O(_0075_)
  );
INV  _0895_ (
    .I(RSTn),
    .O(_0076_)
  );
INV  _0896_ (
    .I(RSTn),
    .O(_0077_)
  );
INV  _0897_ (
    .I(RSTn),
    .O(_0078_)
  );
INV  _0898_ (
    .I(RSTn),
    .O(_0079_)
  );
INV  _0899_ (
    .I(RSTn),
    .O(_0080_)
  );
INV  _0900_ (
    .I(RSTn),
    .O(_0081_)
  );
INV  _0901_ (
    .I(RSTn),
    .O(_0082_)
  );
INV  _0902_ (
    .I(RSTn),
    .O(_0083_)
  );
INV  _0903_ (
    .I(RSTn),
    .O(_0084_)
  );
INV  _0904_ (
    .I(RSTn),
    .O(_0085_)
  );
INV  _0905_ (
    .I(RSTn),
    .O(_0086_)
  );
INV  _0906_ (
    .I(RSTn),
    .O(_0087_)
  );
INV  _0907_ (
    .I(RSTn),
    .O(_0088_)
  );
INV  _0908_ (
    .I(RSTn),
    .O(_0089_)
  );
INV  _0909_ (
    .I(RSTn),
    .O(_0090_)
  );
INV  _0910_ (
    .I(RSTn),
    .O(_0091_)
  );
INV  _0911_ (
    .I(RSTn),
    .O(_0092_)
  );
INV  _0912_ (
    .I(RSTn),
    .O(_0093_)
  );
INV  _0913_ (
    .I(RSTn),
    .O(_0094_)
  );
INV  _0914_ (
    .I(RSTn),
    .O(_0095_)
  );
INV  _0915_ (
    .I(RSTn),
    .O(_0096_)
  );
INV  _0916_ (
    .I(RSTn),
    .O(_0097_)
  );
INV  _0917_ (
    .I(RSTn),
    .O(_0098_)
  );
INV  _0918_ (
    .I(RSTn),
    .O(_0099_)
  );
INV  _0919_ (
    .I(RSTn),
    .O(_0100_)
  );
INV  _0920_ (
    .I(RSTn),
    .O(_0101_)
  );
INV  _0921_ (
    .I(RSTn),
    .O(_0102_)
  );
INV  _0922_ (
    .I(RSTn),
    .O(_0103_)
  );
INV  _0923_ (
    .I(RSTn),
    .O(_0104_)
  );
INV  _0924_ (
    .I(RSTn),
    .O(_0105_)
  );
INV  _0925_ (
    .I(RSTn),
    .O(_0106_)
  );
INV  _0926_ (
    .I(RSTn),
    .O(_0107_)
  );
INV  _0927_ (
    .I(RSTn),
    .O(_0108_)
  );
INV  _0928_ (
    .I(RSTn),
    .O(_0109_)
  );
INV  _0929_ (
    .I(RSTn),
    .O(_0110_)
  );
INV  _0930_ (
    .I(RSTn),
    .O(_0111_)
  );
INV  _0931_ (
    .I(RSTn),
    .O(_0112_)
  );
INV  _0932_ (
    .I(RSTn),
    .O(_0113_)
  );
INV  _0933_ (
    .I(RSTn),
    .O(_0114_)
  );
INV  _0934_ (
    .I(RSTn),
    .O(_0115_)
  );
INV  _0935_ (
    .I(RSTn),
    .O(_0116_)
  );
INV  _0936_ (
    .I(RSTn),
    .O(_0117_)
  );
INV  _0937_ (
    .I(RSTn),
    .O(_0118_)
  );
INV  _0938_ (
    .I(RSTn),
    .O(_0119_)
  );
INV  _0939_ (
    .I(RSTn),
    .O(_0120_)
  );
INV  _0940_ (
    .I(RSTn),
    .O(_0121_)
  );
INV  _0941_ (
    .I(RSTn),
    .O(_0122_)
  );
INV  _0942_ (
    .I(RSTn),
    .O(_0123_)
  );
INV  _0943_ (
    .I(RSTn),
    .O(_0124_)
  );
INV  _0944_ (
    .I(RSTn),
    .O(_0125_)
  );
INV  _0945_ (
    .I(RSTn),
    .O(_0126_)
  );
INV  _0946_ (
    .I(RSTn),
    .O(_0127_)
  );
INV  _0947_ (
    .I(RSTn),
    .O(_0128_)
  );
INV  _0948_ (
    .I(RSTn),
    .O(_0129_)
  );
INV  _0949_ (
    .I(RSTn),
    .O(_0130_)
  );
INV  _0950_ (
    .I(RSTn),
    .O(_0131_)
  );
INV  _0951_ (
    .I(RSTn),
    .O(_0132_)
  );
INV  _0952_ (
    .I(RSTn),
    .O(_0133_)
  );
INV  _0953_ (
    .I(RSTn),
    .O(_0134_)
  );
INV  _0954_ (
    .I(RSTn),
    .O(_0135_)
  );
INV  _0955_ (
    .I(RSTn),
    .O(_0136_)
  );
INV  _0956_ (
    .I(RSTn),
    .O(_0137_)
  );
INV  _0957_ (
    .I(RSTn),
    .O(_0138_)
  );
INV  _0958_ (
    .I(RSTn),
    .O(_0139_)
  );
INV  _0959_ (
    .I(RSTn),
    .O(_0140_)
  );
INV  _0960_ (
    .I(RSTn),
    .O(_0141_)
  );
INV  _0961_ (
    .I(RSTn),
    .O(_0142_)
  );
INV  _0962_ (
    .I(RSTn),
    .O(_0143_)
  );
INV  _0963_ (
    .I(RSTn),
    .O(_0144_)
  );
INV  _0964_ (
    .I(RSTn),
    .O(_0145_)
  );
INV  _0965_ (
    .I(RSTn),
    .O(_0146_)
  );
INV  _0966_ (
    .I(RSTn),
    .O(_0147_)
  );
INV  _0967_ (
    .I(RSTn),
    .O(_0148_)
  );
INV  _0968_ (
    .I(RSTn),
    .O(_0149_)
  );
INV  _0969_ (
    .I(RSTn),
    .O(_0150_)
  );
INV  _0970_ (
    .I(RSTn),
    .O(_0151_)
  );
INV  _0971_ (
    .I(RSTn),
    .O(_0152_)
  );
INV  _0972_ (
    .I(RSTn),
    .O(_0153_)
  );
INV  _0973_ (
    .I(RSTn),
    .O(_0154_)
  );
INV  _0974_ (
    .I(RSTn),
    .O(_0155_)
  );
INV  _0975_ (
    .I(RSTn),
    .O(_0156_)
  );
INV  _0976_ (
    .I(RSTn),
    .O(_0157_)
  );
INV  _0977_ (
    .I(RSTn),
    .O(_0158_)
  );
INV  _0978_ (
    .I(RSTn),
    .O(_0159_)
  );
INV  _0979_ (
    .I(RSTn),
    .O(_0160_)
  );
INV  _0980_ (
    .I(RSTn),
    .O(_0161_)
  );
INV  _0981_ (
    .I(RSTn),
    .O(_0162_)
  );
INV  _0982_ (
    .I(RSTn),
    .O(_0163_)
  );
INV  _0983_ (
    .I(RSTn),
    .O(_0164_)
  );
INV  _0984_ (
    .I(RSTn),
    .O(_0165_)
  );
INV  _0985_ (
    .I(RSTn),
    .O(_0166_)
  );
INV  _0986_ (
    .I(RSTn),
    .O(_0167_)
  );
INV  _0987_ (
    .I(RSTn),
    .O(_0168_)
  );
INV  _0988_ (
    .I(RSTn),
    .O(_0169_)
  );
INV  _0989_ (
    .I(RSTn),
    .O(_0170_)
  );
INV  _0990_ (
    .I(RSTn),
    .O(_0171_)
  );
INV  _0991_ (
    .I(RSTn),
    .O(_0172_)
  );
INV  _0992_ (
    .I(RSTn),
    .O(_0173_)
  );
INV  _0993_ (
    .I(RSTn),
    .O(_0174_)
  );
INV  _0994_ (
    .I(RSTn),
    .O(_0175_)
  );
INV  _0995_ (
    .I(RSTn),
    .O(_0176_)
  );
INV  _0996_ (
    .I(RSTn),
    .O(_0177_)
  );
INV  _0997_ (
    .I(RSTn),
    .O(_0178_)
  );
INV  _0998_ (
    .I(RSTn),
    .O(_0179_)
  );
INV  _0999_ (
    .I(RSTn),
    .O(_0180_)
  );
INV  _1000_ (
    .I(RSTn),
    .O(_0181_)
  );
INV  _1001_ (
    .I(RSTn),
    .O(_0182_)
  );
INV  _1002_ (
    .I(RSTn),
    .O(_0183_)
  );
INV  _1003_ (
    .I(RSTn),
    .O(_0184_)
  );
INV  _1004_ (
    .I(RSTn),
    .O(_0185_)
  );
INV  _1005_ (
    .I(RSTn),
    .O(_0186_)
  );
INV  _1006_ (
    .I(RSTn),
    .O(_0187_)
  );
INV  _1007_ (
    .I(RSTn),
    .O(_0188_)
  );
INV  _1008_ (
    .I(RSTn),
    .O(_0189_)
  );
INV  _1009_ (
    .I(RSTn),
    .O(_0190_)
  );
INV  _1010_ (
    .I(RSTn),
    .O(_0191_)
  );
INV  _1011_ (
    .I(RSTn),
    .O(_0192_)
  );
INV  _1012_ (
    .I(RSTn),
    .O(_0193_)
  );
INV  _1013_ (
    .I(RSTn),
    .O(_0194_)
  );
INV  _1014_ (
    .I(RSTn),
    .O(_0195_)
  );
INV  _1015_ (
    .I(RSTn),
    .O(_0196_)
  );
INV  _1016_ (
    .I(RSTn),
    .O(_0197_)
  );
INV  _1017_ (
    .I(RSTn),
    .O(_0198_)
  );
INV  _1018_ (
    .I(RSTn),
    .O(_0199_)
  );
INV  _1019_ (
    .I(RSTn),
    .O(_0200_)
  );
INV  _1020_ (
    .I(RSTn),
    .O(_0201_)
  );
INV  _1021_ (
    .I(RSTn),
    .O(_0202_)
  );
INV  _1022_ (
    .I(RSTn),
    .O(_0203_)
  );
INV  _1023_ (
    .I(RSTn),
    .O(_0204_)
  );
INV  _1024_ (
    .I(RSTn),
    .O(_0205_)
  );
INV  _1025_ (
    .I(RSTn),
    .O(_0206_)
  );
INV  _1026_ (
    .I(RSTn),
    .O(_0207_)
  );
INV  _1027_ (
    .I(RSTn),
    .O(_0208_)
  );
INV  _1028_ (
    .I(RSTn),
    .O(_0209_)
  );
INV  _1029_ (
    .I(RSTn),
    .O(_0210_)
  );
INV  _1030_ (
    .I(RSTn),
    .O(_0211_)
  );
INV  _1031_ (
    .I(RSTn),
    .O(_0212_)
  );
INV  _1032_ (
    .I(RSTn),
    .O(_0213_)
  );
INV  _1033_ (
    .I(RSTn),
    .O(_0214_)
  );
INV  _1034_ (
    .I(RSTn),
    .O(_0215_)
  );
INV  _1035_ (
    .I(RSTn),
    .O(_0216_)
  );
INV  _1036_ (
    .I(RSTn),
    .O(_0217_)
  );
INV  _1037_ (
    .I(RSTn),
    .O(_0218_)
  );
INV  _1038_ (
    .I(RSTn),
    .O(_0219_)
  );
INV  _1039_ (
    .I(RSTn),
    .O(_0220_)
  );
INV  _1040_ (
    .I(RSTn),
    .O(_0221_)
  );
INV  _1041_ (
    .I(RSTn),
    .O(_0222_)
  );
INV  _1042_ (
    .I(RSTn),
    .O(_0223_)
  );
INV  _1043_ (
    .I(RSTn),
    .O(_0224_)
  );
INV  _1044_ (
    .I(RSTn),
    .O(_0225_)
  );
INV  _1045_ (
    .I(RSTn),
    .O(_0226_)
  );
INV  _1046_ (
    .I(RSTn),
    .O(_0227_)
  );
INV  _1047_ (
    .I(RSTn),
    .O(_0228_)
  );
INV  _1048_ (
    .I(RSTn),
    .O(_0229_)
  );
INV  _1049_ (
    .I(RSTn),
    .O(_0230_)
  );
INV  _1050_ (
    .I(RSTn),
    .O(_0231_)
  );
INV  _1051_ (
    .I(RSTn),
    .O(_0232_)
  );
INV  _1052_ (
    .I(RSTn),
    .O(_0233_)
  );
INV  _1053_ (
    .I(RSTn),
    .O(_0234_)
  );
INV  _1054_ (
    .I(RSTn),
    .O(_0235_)
  );
INV  _1055_ (
    .I(RSTn),
    .O(_0236_)
  );
INV  _1056_ (
    .I(RSTn),
    .O(_0237_)
  );
INV  _1057_ (
    .I(RSTn),
    .O(_0238_)
  );
INV  _1058_ (
    .I(RSTn),
    .O(_0239_)
  );
INV  _1059_ (
    .I(RSTn),
    .O(_0240_)
  );
INV  _1060_ (
    .I(RSTn),
    .O(_0241_)
  );
INV  _1061_ (
    .I(RSTn),
    .O(_0242_)
  );
INV  _1062_ (
    .I(RSTn),
    .O(_0243_)
  );
INV  _1063_ (
    .I(RSTn),
    .O(_0244_)
  );
INV  _1064_ (
    .I(RSTn),
    .O(_0245_)
  );
INV  _1065_ (
    .I(RSTn),
    .O(_0246_)
  );
INV  _1066_ (
    .I(RSTn),
    .O(_0247_)
  );
INV  _1067_ (
    .I(RSTn),
    .O(_0248_)
  );
INV  _1068_ (
    .I(RSTn),
    .O(_0249_)
  );
INV  _1069_ (
    .I(RSTn),
    .O(_0250_)
  );
INV  _1070_ (
    .I(RSTn),
    .O(_0251_)
  );
INV  _1071_ (
    .I(RSTn),
    .O(_0252_)
  );
INV  _1072_ (
    .I(RSTn),
    .O(_0253_)
  );
INV  _1073_ (
    .I(RSTn),
    .O(_0254_)
  );
INV  _1074_ (
    .I(RSTn),
    .O(_0255_)
  );
INV  _1075_ (
    .I(RSTn),
    .O(_0256_)
  );
INV  _1076_ (
    .I(RSTn),
    .O(_0257_)
  );
INV  _1077_ (
    .I(RSTn),
    .O(_0258_)
  );
INV  _1078_ (
    .I(RSTn),
    .O(_0259_)
  );
INV  _1079_ (
    .I(RSTn),
    .O(_0260_)
  );
INV  _1080_ (
    .I(RSTn),
    .O(_0261_)
  );
INV  _1081_ (
    .I(RSTn),
    .O(_0262_)
  );
INV  _1082_ (
    .I(RSTn),
    .O(_0263_)
  );
INV  _1083_ (
    .I(RSTn),
    .O(_0264_)
  );
INV  _1084_ (
    .I(RSTn),
    .O(_0265_)
  );
INV  _1085_ (
    .I(RSTn),
    .O(_0266_)
  );
INV  _1086_ (
    .I(RSTn),
    .O(_0267_)
  );
INV  _1087_ (
    .I(RSTn),
    .O(_0268_)
  );
INV  _1088_ (
    .I(RSTn),
    .O(_0269_)
  );
INV  _1089_ (
    .I(RSTn),
    .O(_0270_)
  );
INV  _1090_ (
    .I(RSTn),
    .O(_0271_)
  );
INV  _1091_ (
    .I(RSTn),
    .O(_0272_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1092_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0403_),
    .Q(Drg[0]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1093_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0442_),
    .Q(Drg[1]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1094_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0453_),
    .Q(Drg[2]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1095_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0464_),
    .Q(Drg[3]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1096_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0475_),
    .Q(Drg[4]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1097_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0486_),
    .Q(Drg[5]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1098_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0497_),
    .Q(Drg[6]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1099_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0508_),
    .Q(Drg[7]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1100_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0519_),
    .Q(Drg[8]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1101_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0530_),
    .Q(Drg[9]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1102_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0414_),
    .Q(Drg[10]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1103_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0425_),
    .Q(Drg[11]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1104_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0434_),
    .Q(Drg[12]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1105_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0435_),
    .Q(Drg[13]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1106_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0436_),
    .Q(Drg[14]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1107_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0437_),
    .Q(Drg[15]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1108_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0438_),
    .Q(Drg[16]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1109_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0439_),
    .Q(Drg[17]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1110_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0440_),
    .Q(Drg[18]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1111_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0441_),
    .Q(Drg[19]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1112_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0443_),
    .Q(Drg[20]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1113_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0444_),
    .Q(Drg[21]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1114_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0445_),
    .Q(Drg[22]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1115_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0446_),
    .Q(Drg[23]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1116_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0447_),
    .Q(Drg[24]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1117_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0448_),
    .Q(Drg[25]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1118_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0449_),
    .Q(Drg[26]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1119_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0450_),
    .Q(Drg[27]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1120_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0451_),
    .Q(Drg[28]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1121_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0452_),
    .Q(Drg[29]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1122_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0454_),
    .Q(Drg[30]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1123_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0455_),
    .Q(Drg[31]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1124_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0456_),
    .Q(Drg[32]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1125_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0457_),
    .Q(Drg[33]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1126_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0458_),
    .Q(Drg[34]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1127_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0459_),
    .Q(Drg[35]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1128_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0460_),
    .Q(Drg[36]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1129_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0461_),
    .Q(Drg[37]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1130_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0462_),
    .Q(Drg[38]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1131_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0463_),
    .Q(Drg[39]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1132_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0465_),
    .Q(Drg[40]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1133_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0466_),
    .Q(Drg[41]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1134_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0467_),
    .Q(Drg[42]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1135_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0468_),
    .Q(Drg[43]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1136_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0469_),
    .Q(Drg[44]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1137_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0470_),
    .Q(Drg[45]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1138_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0471_),
    .Q(Drg[46]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1139_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0472_),
    .Q(Drg[47]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1140_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0473_),
    .Q(Drg[48]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1141_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0474_),
    .Q(Drg[49]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1142_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0476_),
    .Q(Drg[50]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1143_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0477_),
    .Q(Drg[51]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1144_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0478_),
    .Q(Drg[52]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1145_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0479_),
    .Q(Drg[53]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1146_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0480_),
    .Q(Drg[54]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1147_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0481_),
    .Q(Drg[55]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1148_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0482_),
    .Q(Drg[56]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1149_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0483_),
    .Q(Drg[57]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1150_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0484_),
    .Q(Drg[58]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1151_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0485_),
    .Q(Drg[59]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1152_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0487_),
    .Q(Drg[60]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1153_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0488_),
    .Q(Drg[61]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1154_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0489_),
    .Q(Drg[62]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1155_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0490_),
    .Q(Drg[63]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1156_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0491_),
    .Q(Drg[64]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1157_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0492_),
    .Q(Drg[65]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1158_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0493_),
    .Q(Drg[66]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1159_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0494_),
    .Q(Drg[67]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1160_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0495_),
    .Q(Drg[68]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1161_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0496_),
    .Q(Drg[69]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1162_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0498_),
    .Q(Drg[70]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1163_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0499_),
    .Q(Drg[71]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1164_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0500_),
    .Q(Drg[72]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1165_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0501_),
    .Q(Drg[73]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1166_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0502_),
    .Q(Drg[74]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1167_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0503_),
    .Q(Drg[75]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1168_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0504_),
    .Q(Drg[76]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1169_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0505_),
    .Q(Drg[77]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1170_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0506_),
    .Q(Drg[78]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1171_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0507_),
    .Q(Drg[79]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1172_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0509_),
    .Q(Drg[80]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1173_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0510_),
    .Q(Drg[81]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1174_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0511_),
    .Q(Drg[82]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1175_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0512_),
    .Q(Drg[83]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1176_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0513_),
    .Q(Drg[84]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1177_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0514_),
    .Q(Drg[85]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1178_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0515_),
    .Q(Drg[86]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1179_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0516_),
    .Q(Drg[87]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1180_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0517_),
    .Q(Drg[88]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1181_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0518_),
    .Q(Drg[89]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1182_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0520_),
    .Q(Drg[90]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1183_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0521_),
    .Q(Drg[91]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1184_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0522_),
    .Q(Drg[92]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1185_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0523_),
    .Q(Drg[93]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1186_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0524_),
    .Q(Drg[94]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1187_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0525_),
    .Q(Drg[95]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1188_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0526_),
    .Q(Drg[96]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1189_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0527_),
    .Q(Drg[97]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1190_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0528_),
    .Q(Drg[98]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1191_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0529_),
    .Q(Drg[99]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1192_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0404_),
    .Q(Drg[100]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1193_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0405_),
    .Q(Drg[101]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1194_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0406_),
    .Q(Drg[102]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1195_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0407_),
    .Q(Drg[103]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1196_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0408_),
    .Q(Drg[104]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1197_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0409_),
    .Q(Drg[105]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1198_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0410_),
    .Q(Drg[106]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1199_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0411_),
    .Q(Drg[107]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1200_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0412_),
    .Q(Drg[108]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1201_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0413_),
    .Q(Drg[109]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1202_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0415_),
    .Q(Drg[110]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1203_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0416_),
    .Q(Drg[111]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1204_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0417_),
    .Q(Drg[112]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1205_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0418_),
    .Q(Drg[113]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1206_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0419_),
    .Q(Drg[114]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1207_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0420_),
    .Q(Drg[115]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1208_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0421_),
    .Q(Drg[116]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1209_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0422_),
    .Q(Drg[117]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1210_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0423_),
    .Q(Drg[118]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1211_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0424_),
    .Q(Drg[119]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1212_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0426_),
    .Q(Drg[120]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1213_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0427_),
    .Q(Drg[121]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1214_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0428_),
    .Q(Drg[122]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1215_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0429_),
    .Q(Drg[123]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1216_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0430_),
    .Q(Drg[124]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1217_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0431_),
    .Q(Drg[125]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1218_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0432_),
    .Q(Drg[126]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1219_ (
    .C(CLK),
    .CE(_0010_),
    .D(_0433_),
    .Q(Drg[127]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1220_ (
    .C(CLK),
    .CE(_0012_),
    .D(_0531_),
    .Q(Rrg[0]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1221_ (
    .C(CLK),
    .CE(_0012_),
    .D(_0532_),
    .Q(Rrg[1]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1222_ (
    .C(CLK),
    .CE(_0012_),
    .D(_0533_),
    .Q(Rrg[2]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1223_ (
    .C(CLK),
    .CE(_0012_),
    .D(_0534_),
    .Q(Rrg[3]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1224_ (
    .C(CLK),
    .CE(_0012_),
    .D(_0535_),
    .Q(Rrg[4]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1225_ (
    .C(CLK),
    .CE(_0012_),
    .D(_0536_),
    .Q(Rrg[5]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1226_ (
    .C(CLK),
    .CE(_0012_),
    .D(_0537_),
    .Q(Rrg[6]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1227_ (
    .C(CLK),
    .CE(_0012_),
    .D(_0538_),
    .Q(Rrg[7]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1228_ (
    .C(CLK),
    .CE(_0012_),
    .D(_0539_),
    .Q(Rrg[8]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1229_ (
    .C(CLK),
    .CE(_0011_),
    .D(_0540_),
    .Q(Rrg[9]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1230_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[0]),
    .Q(Krg[0]),
    .R(_0014_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1231_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[1]),
    .Q(Krg[1]),
    .R(_0015_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1232_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[2]),
    .Q(Krg[2]),
    .R(_0016_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1233_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[3]),
    .Q(Krg[3]),
    .R(_0017_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1234_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[4]),
    .Q(Krg[4]),
    .R(_0018_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1235_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[5]),
    .Q(Krg[5]),
    .R(_0019_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1236_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[6]),
    .Q(Krg[6]),
    .R(_0020_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1237_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[7]),
    .Q(Krg[7]),
    .R(_0021_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1238_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[8]),
    .Q(Krg[8]),
    .R(_0022_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1239_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[9]),
    .Q(Krg[9]),
    .R(_0023_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1240_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[10]),
    .Q(Krg[10]),
    .R(_0024_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1241_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[11]),
    .Q(Krg[11]),
    .R(_0025_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1242_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[12]),
    .Q(Krg[12]),
    .R(_0026_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1243_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[13]),
    .Q(Krg[13]),
    .R(_0027_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1244_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[14]),
    .Q(Krg[14]),
    .R(_0028_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1245_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[15]),
    .Q(Krg[15]),
    .R(_0029_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1246_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[16]),
    .Q(Krg[16]),
    .R(_0030_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1247_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[17]),
    .Q(Krg[17]),
    .R(_0031_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1248_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[18]),
    .Q(Krg[18]),
    .R(_0032_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1249_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[19]),
    .Q(Krg[19]),
    .R(_0033_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1250_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[20]),
    .Q(Krg[20]),
    .R(_0034_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1251_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[21]),
    .Q(Krg[21]),
    .R(_0035_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1252_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[22]),
    .Q(Krg[22]),
    .R(_0036_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1253_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[23]),
    .Q(Krg[23]),
    .R(_0037_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1254_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[24]),
    .Q(Krg[24]),
    .R(_0038_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1255_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[25]),
    .Q(Krg[25]),
    .R(_0039_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1256_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[26]),
    .Q(Krg[26]),
    .R(_0040_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1257_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[27]),
    .Q(Krg[27]),
    .R(_0041_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1258_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[28]),
    .Q(Krg[28]),
    .R(_0042_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1259_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[29]),
    .Q(Krg[29]),
    .R(_0043_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1260_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[30]),
    .Q(Krg[30]),
    .R(_0044_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1261_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[31]),
    .Q(Krg[31]),
    .R(_0045_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1262_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[32]),
    .Q(Krg[32]),
    .R(_0046_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1263_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[33]),
    .Q(Krg[33]),
    .R(_0047_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1264_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[34]),
    .Q(Krg[34]),
    .R(_0048_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1265_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[35]),
    .Q(Krg[35]),
    .R(_0049_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1266_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[36]),
    .Q(Krg[36]),
    .R(_0050_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1267_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[37]),
    .Q(Krg[37]),
    .R(_0051_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1268_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[38]),
    .Q(Krg[38]),
    .R(_0052_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1269_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[39]),
    .Q(Krg[39]),
    .R(_0053_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1270_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[40]),
    .Q(Krg[40]),
    .R(_0054_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1271_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[41]),
    .Q(Krg[41]),
    .R(_0055_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1272_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[42]),
    .Q(Krg[42]),
    .R(_0056_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1273_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[43]),
    .Q(Krg[43]),
    .R(_0057_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1274_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[44]),
    .Q(Krg[44]),
    .R(_0058_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1275_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[45]),
    .Q(Krg[45]),
    .R(_0059_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1276_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[46]),
    .Q(Krg[46]),
    .R(_0060_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1277_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[47]),
    .Q(Krg[47]),
    .R(_0061_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1278_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[48]),
    .Q(Krg[48]),
    .R(_0062_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1279_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[49]),
    .Q(Krg[49]),
    .R(_0063_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1280_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[50]),
    .Q(Krg[50]),
    .R(_0064_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1281_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[51]),
    .Q(Krg[51]),
    .R(_0065_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1282_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[52]),
    .Q(Krg[52]),
    .R(_0066_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1283_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[53]),
    .Q(Krg[53]),
    .R(_0067_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1284_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[54]),
    .Q(Krg[54]),
    .R(_0068_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1285_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[55]),
    .Q(Krg[55]),
    .R(_0069_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1286_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[56]),
    .Q(Krg[56]),
    .R(_0070_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1287_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[57]),
    .Q(Krg[57]),
    .R(_0071_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1288_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[58]),
    .Q(Krg[58]),
    .R(_0072_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1289_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[59]),
    .Q(Krg[59]),
    .R(_0073_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1290_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[60]),
    .Q(Krg[60]),
    .R(_0074_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1291_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[61]),
    .Q(Krg[61]),
    .R(_0075_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1292_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[62]),
    .Q(Krg[62]),
    .R(_0076_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1293_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[63]),
    .Q(Krg[63]),
    .R(_0077_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1294_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[64]),
    .Q(Krg[64]),
    .R(_0078_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1295_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[65]),
    .Q(Krg[65]),
    .R(_0079_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1296_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[66]),
    .Q(Krg[66]),
    .R(_0080_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1297_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[67]),
    .Q(Krg[67]),
    .R(_0081_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1298_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[68]),
    .Q(Krg[68]),
    .R(_0082_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1299_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[69]),
    .Q(Krg[69]),
    .R(_0083_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1300_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[70]),
    .Q(Krg[70]),
    .R(_0084_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1301_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[71]),
    .Q(Krg[71]),
    .R(_0085_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1302_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[72]),
    .Q(Krg[72]),
    .R(_0086_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1303_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[73]),
    .Q(Krg[73]),
    .R(_0087_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1304_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[74]),
    .Q(Krg[74]),
    .R(_0088_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1305_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[75]),
    .Q(Krg[75]),
    .R(_0089_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1306_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[76]),
    .Q(Krg[76]),
    .R(_0090_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1307_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[77]),
    .Q(Krg[77]),
    .R(_0091_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1308_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[78]),
    .Q(Krg[78]),
    .R(_0092_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1309_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[79]),
    .Q(Krg[79]),
    .R(_0093_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1310_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[80]),
    .Q(Krg[80]),
    .R(_0094_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1311_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[81]),
    .Q(Krg[81]),
    .R(_0095_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1312_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[82]),
    .Q(Krg[82]),
    .R(_0096_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1313_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[83]),
    .Q(Krg[83]),
    .R(_0097_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1314_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[84]),
    .Q(Krg[84]),
    .R(_0098_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1315_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[85]),
    .Q(Krg[85]),
    .R(_0099_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1316_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[86]),
    .Q(Krg[86]),
    .R(_0100_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1317_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[87]),
    .Q(Krg[87]),
    .R(_0101_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1318_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[88]),
    .Q(Krg[88]),
    .R(_0102_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1319_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[89]),
    .Q(Krg[89]),
    .R(_0103_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1320_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[90]),
    .Q(Krg[90]),
    .R(_0104_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1321_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[91]),
    .Q(Krg[91]),
    .R(_0105_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1322_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[92]),
    .Q(Krg[92]),
    .R(_0106_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1323_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[93]),
    .Q(Krg[93]),
    .R(_0107_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1324_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[94]),
    .Q(Krg[94]),
    .R(_0108_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1325_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[95]),
    .Q(Krg[95]),
    .R(_0109_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1326_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[96]),
    .Q(Krg[96]),
    .R(_0110_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1327_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[97]),
    .Q(Krg[97]),
    .R(_0111_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1328_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[98]),
    .Q(Krg[98]),
    .R(_0112_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1329_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[99]),
    .Q(Krg[99]),
    .R(_0113_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1330_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[100]),
    .Q(Krg[100]),
    .R(_0114_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1331_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[101]),
    .Q(Krg[101]),
    .R(_0115_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1332_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[102]),
    .Q(Krg[102]),
    .R(_0116_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1333_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[103]),
    .Q(Krg[103]),
    .R(_0117_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1334_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[104]),
    .Q(Krg[104]),
    .R(_0118_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1335_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[105]),
    .Q(Krg[105]),
    .R(_0119_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1336_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[106]),
    .Q(Krg[106]),
    .R(_0120_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1337_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[107]),
    .Q(Krg[107]),
    .R(_0121_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1338_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[108]),
    .Q(Krg[108]),
    .R(_0122_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1339_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[109]),
    .Q(Krg[109]),
    .R(_0123_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1340_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[110]),
    .Q(Krg[110]),
    .R(_0124_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1341_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[111]),
    .Q(Krg[111]),
    .R(_0125_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1342_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[112]),
    .Q(Krg[112]),
    .R(_0126_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1343_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[113]),
    .Q(Krg[113]),
    .R(_0127_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1344_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[114]),
    .Q(Krg[114]),
    .R(_0128_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1345_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[115]),
    .Q(Krg[115]),
    .R(_0129_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1346_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[116]),
    .Q(Krg[116]),
    .R(_0130_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1347_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[117]),
    .Q(Krg[117]),
    .R(_0131_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1348_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[118]),
    .Q(Krg[118]),
    .R(_0132_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1349_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[119]),
    .Q(Krg[119]),
    .R(_0133_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1350_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[120]),
    .Q(Krg[120]),
    .R(_0134_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1351_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[121]),
    .Q(Krg[121]),
    .R(_0135_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1352_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[122]),
    .Q(Krg[122]),
    .R(_0136_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1353_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[123]),
    .Q(Krg[123]),
    .R(_0137_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1354_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[124]),
    .Q(Krg[124]),
    .R(_0138_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1355_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[125]),
    .Q(Krg[125]),
    .R(_0139_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1356_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[126]),
    .Q(Krg[126]),
    .R(_0140_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1357_ (
    .C(CLK),
    .CE(_0009_),
    .D(KrgX[127]),
    .Q(Krg[127]),
    .R(_0141_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1358_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0275_),
    .Q(KrgX[0]),
    .R(_0142_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1359_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0314_),
    .Q(KrgX[1]),
    .R(_0143_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1360_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0325_),
    .Q(KrgX[2]),
    .R(_0144_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1361_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0336_),
    .Q(KrgX[3]),
    .R(_0145_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1362_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0347_),
    .Q(KrgX[4]),
    .R(_0146_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1363_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0358_),
    .Q(KrgX[5]),
    .R(_0147_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1364_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0369_),
    .Q(KrgX[6]),
    .R(_0148_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1365_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0380_),
    .Q(KrgX[7]),
    .R(_0149_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1366_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0391_),
    .Q(KrgX[8]),
    .R(_0150_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1367_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0402_),
    .Q(KrgX[9]),
    .R(_0151_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1368_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0286_),
    .Q(KrgX[10]),
    .R(_0152_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1369_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0297_),
    .Q(KrgX[11]),
    .R(_0153_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1370_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0306_),
    .Q(KrgX[12]),
    .R(_0154_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1371_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0307_),
    .Q(KrgX[13]),
    .R(_0155_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1372_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0308_),
    .Q(KrgX[14]),
    .R(_0156_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1373_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0309_),
    .Q(KrgX[15]),
    .R(_0157_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1374_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0310_),
    .Q(KrgX[16]),
    .R(_0158_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1375_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0311_),
    .Q(KrgX[17]),
    .R(_0159_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1376_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0312_),
    .Q(KrgX[18]),
    .R(_0160_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1377_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0313_),
    .Q(KrgX[19]),
    .R(_0161_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1378_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0315_),
    .Q(KrgX[20]),
    .R(_0162_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1379_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0316_),
    .Q(KrgX[21]),
    .R(_0163_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1380_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0317_),
    .Q(KrgX[22]),
    .R(_0164_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1381_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0318_),
    .Q(KrgX[23]),
    .R(_0165_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1382_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0319_),
    .Q(KrgX[24]),
    .R(_0166_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1383_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0320_),
    .Q(KrgX[25]),
    .R(_0167_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1384_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0321_),
    .Q(KrgX[26]),
    .R(_0168_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1385_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0322_),
    .Q(KrgX[27]),
    .R(_0169_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1386_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0323_),
    .Q(KrgX[28]),
    .R(_0170_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1387_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0324_),
    .Q(KrgX[29]),
    .R(_0171_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1388_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0326_),
    .Q(KrgX[30]),
    .R(_0172_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1389_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0327_),
    .Q(KrgX[31]),
    .R(_0173_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1390_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0328_),
    .Q(KrgX[32]),
    .R(_0174_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1391_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0329_),
    .Q(KrgX[33]),
    .R(_0175_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1392_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0330_),
    .Q(KrgX[34]),
    .R(_0176_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1393_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0331_),
    .Q(KrgX[35]),
    .R(_0177_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1394_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0332_),
    .Q(KrgX[36]),
    .R(_0178_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1395_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0333_),
    .Q(KrgX[37]),
    .R(_0179_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1396_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0334_),
    .Q(KrgX[38]),
    .R(_0180_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1397_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0335_),
    .Q(KrgX[39]),
    .R(_0181_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1398_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0337_),
    .Q(KrgX[40]),
    .R(_0182_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1399_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0338_),
    .Q(KrgX[41]),
    .R(_0183_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1400_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0339_),
    .Q(KrgX[42]),
    .R(_0184_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1401_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0340_),
    .Q(KrgX[43]),
    .R(_0185_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1402_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0341_),
    .Q(KrgX[44]),
    .R(_0186_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1403_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0342_),
    .Q(KrgX[45]),
    .R(_0187_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1404_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0343_),
    .Q(KrgX[46]),
    .R(_0188_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1405_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0344_),
    .Q(KrgX[47]),
    .R(_0189_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1406_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0345_),
    .Q(KrgX[48]),
    .R(_0190_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1407_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0346_),
    .Q(KrgX[49]),
    .R(_0191_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1408_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0348_),
    .Q(KrgX[50]),
    .R(_0192_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1409_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0349_),
    .Q(KrgX[51]),
    .R(_0193_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1410_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0350_),
    .Q(KrgX[52]),
    .R(_0194_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1411_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0351_),
    .Q(KrgX[53]),
    .R(_0195_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1412_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0352_),
    .Q(KrgX[54]),
    .R(_0196_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1413_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0353_),
    .Q(KrgX[55]),
    .R(_0197_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1414_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0354_),
    .Q(KrgX[56]),
    .R(_0198_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1415_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0355_),
    .Q(KrgX[57]),
    .R(_0199_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1416_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0356_),
    .Q(KrgX[58]),
    .R(_0200_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1417_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0357_),
    .Q(KrgX[59]),
    .R(_0201_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1418_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0359_),
    .Q(KrgX[60]),
    .R(_0202_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1419_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0360_),
    .Q(KrgX[61]),
    .R(_0203_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1420_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0361_),
    .Q(KrgX[62]),
    .R(_0204_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1421_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0362_),
    .Q(KrgX[63]),
    .R(_0205_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1422_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0363_),
    .Q(KrgX[64]),
    .R(_0206_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1423_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0364_),
    .Q(KrgX[65]),
    .R(_0207_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1424_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0365_),
    .Q(KrgX[66]),
    .R(_0208_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1425_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0366_),
    .Q(KrgX[67]),
    .R(_0209_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1426_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0367_),
    .Q(KrgX[68]),
    .R(_0210_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1427_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0368_),
    .Q(KrgX[69]),
    .R(_0211_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1428_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0370_),
    .Q(KrgX[70]),
    .R(_0212_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1429_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0371_),
    .Q(KrgX[71]),
    .R(_0213_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1430_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0372_),
    .Q(KrgX[72]),
    .R(_0214_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1431_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0373_),
    .Q(KrgX[73]),
    .R(_0215_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1432_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0374_),
    .Q(KrgX[74]),
    .R(_0216_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1433_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0375_),
    .Q(KrgX[75]),
    .R(_0217_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1434_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0376_),
    .Q(KrgX[76]),
    .R(_0218_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1435_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0377_),
    .Q(KrgX[77]),
    .R(_0219_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1436_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0378_),
    .Q(KrgX[78]),
    .R(_0220_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1437_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0379_),
    .Q(KrgX[79]),
    .R(_0221_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1438_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0381_),
    .Q(KrgX[80]),
    .R(_0222_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1439_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0382_),
    .Q(KrgX[81]),
    .R(_0223_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1440_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0383_),
    .Q(KrgX[82]),
    .R(_0224_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1441_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0384_),
    .Q(KrgX[83]),
    .R(_0225_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1442_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0385_),
    .Q(KrgX[84]),
    .R(_0226_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1443_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0386_),
    .Q(KrgX[85]),
    .R(_0227_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1444_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0387_),
    .Q(KrgX[86]),
    .R(_0228_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1445_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0388_),
    .Q(KrgX[87]),
    .R(_0229_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1446_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0389_),
    .Q(KrgX[88]),
    .R(_0230_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1447_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0390_),
    .Q(KrgX[89]),
    .R(_0231_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1448_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0392_),
    .Q(KrgX[90]),
    .R(_0232_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1449_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0393_),
    .Q(KrgX[91]),
    .R(_0233_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1450_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0394_),
    .Q(KrgX[92]),
    .R(_0234_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1451_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0395_),
    .Q(KrgX[93]),
    .R(_0235_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1452_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0396_),
    .Q(KrgX[94]),
    .R(_0236_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1453_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0397_),
    .Q(KrgX[95]),
    .R(_0237_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1454_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0398_),
    .Q(KrgX[96]),
    .R(_0238_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1455_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0399_),
    .Q(KrgX[97]),
    .R(_0239_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1456_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0400_),
    .Q(KrgX[98]),
    .R(_0240_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1457_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0401_),
    .Q(KrgX[99]),
    .R(_0241_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1458_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0276_),
    .Q(KrgX[100]),
    .R(_0242_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1459_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0277_),
    .Q(KrgX[101]),
    .R(_0243_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1460_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0278_),
    .Q(KrgX[102]),
    .R(_0244_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1461_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0279_),
    .Q(KrgX[103]),
    .R(_0245_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1462_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0280_),
    .Q(KrgX[104]),
    .R(_0246_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1463_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0281_),
    .Q(KrgX[105]),
    .R(_0247_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1464_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0282_),
    .Q(KrgX[106]),
    .R(_0248_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1465_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0283_),
    .Q(KrgX[107]),
    .R(_0249_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1466_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0284_),
    .Q(KrgX[108]),
    .R(_0250_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1467_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0285_),
    .Q(KrgX[109]),
    .R(_0251_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1468_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0287_),
    .Q(KrgX[110]),
    .R(_0252_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1469_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0288_),
    .Q(KrgX[111]),
    .R(_0253_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1470_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0289_),
    .Q(KrgX[112]),
    .R(_0254_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1471_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0290_),
    .Q(KrgX[113]),
    .R(_0255_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1472_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0291_),
    .Q(KrgX[114]),
    .R(_0256_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1473_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0292_),
    .Q(KrgX[115]),
    .R(_0257_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1474_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0293_),
    .Q(KrgX[116]),
    .R(_0258_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1475_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0294_),
    .Q(KrgX[117]),
    .R(_0259_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1476_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0295_),
    .Q(KrgX[118]),
    .R(_0260_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1477_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0296_),
    .Q(KrgX[119]),
    .R(_0261_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1478_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0298_),
    .Q(KrgX[120]),
    .R(_0262_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1479_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0299_),
    .Q(KrgX[121]),
    .R(_0263_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1480_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0300_),
    .Q(KrgX[122]),
    .R(_0264_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1481_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0301_),
    .Q(KrgX[123]),
    .R(_0265_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1482_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0302_),
    .Q(KrgX[124]),
    .R(_0266_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1483_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0303_),
    .Q(KrgX[125]),
    .R(_0267_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1484_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0304_),
    .Q(KrgX[126]),
    .R(_0268_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1485_ (
    .C(CLK),
    .CE(_0008_),
    .D(_0305_),
    .Q(KrgX[127]),
    .R(_0269_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1486_ (
    .C(CLK),
    .CE(_0007_),
    .D(_0274_),
    .Q(Kvldrg),
    .R(_0270_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1487_ (
    .C(CLK),
    .CE(_0006_),
    .D(BSYrg),
    .Q(Dvldrg),
    .R(_0271_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _1488_ (
    .C(CLK),
    .CE(EN),
    .D(_0273_),
    .Q(BSYrg),
    .R(_0272_)
  );
AES_Comp_DecCore  DC (
    .Kgen(_0013_),
    .Rrg(Rrg),
    .di(Drg),
    .\do (Dnext),
    .ki(KrgX),
    .ko(Knext)
  );
assign  _0003_[4:0] = { Kvldrg, Rrg[8], _0000_[2:1], Rrg[7] };
assign  { _0541_[5:3], _0541_[1:0] } = { BSYrg, Knext[127], Krdy, Krg[127], Kin[127] };
assign  _0542_[2:0] = { RSTn, _0541_[2], BSYrg };
assign  _0543_[4:1] = { EN, _0000_[1:0], _0000_[2] };
assign  { _0000_[6:5], _0000_[3] } = { BSYrg, Kvldrg, Rrg[9] };
assign  BSY = BSYrg;
assign  Dout = Drg;
assign  Dvld = Dvldrg;
assign  Kvld = Kvldrg;
endmodule
