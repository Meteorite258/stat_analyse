module xS(clk,  in, out);
wire  _000_;
wire  _001_;
wire  _002_;
wire  _003_;
wire  _004_;
wire  _005_;
wire  _006_;
wire  _007_;
wire  _008_;
wire  _009_;
wire  _010_;
wire  _011_;
wire  _012_;
wire  _013_;
wire  _014_;
wire  _015_;
wire  _016_;
wire  _017_;
wire  _018_;
wire  _019_;
wire  _020_;
wire  _021_;
wire  _022_;
wire  _023_;
wire  _024_;
wire  _025_;
wire  _026_;
wire  _027_;
wire  _028_;
wire  _029_;
wire  _030_;
wire  _031_;
wire  _032_;
wire  _033_;
wire  _034_;
wire  _035_;
wire  _036_;
wire  _037_;
wire  _038_;
wire  _039_;
wire  _040_;
wire  _041_;
wire  _042_;
wire  _043_;
wire  _044_;
wire  _045_;
wire  _046_;
wire  _047_;
wire  [7:0] _048_;
input  clk;
input  [7:0] in;
output  [7:0] out;
LUT6  #(
    .INIT(64'h8c9a4ac442f5b9cc)
  ) _049_ (
    .I0(in[0]),
    .I1(in[4]),
    .I2(in[3]),
    .I3(in[7]),
    .I4(in[2]),
    .I5(in[1]),
    .O(_002_)
  );
LUT6  #(
    .INIT(64'h584bd0f93c683d2b)
  ) _050_ (
    .I0(in[0]),
    .I1(in[4]),
    .I2(in[3]),
    .I3(in[7]),
    .I4(in[2]),
    .I5(in[1]),
    .O(_003_)
  );
MUXF7  _051_ (
    .I0(_002_),
    .I1(_003_),
    .O(_000_),
    .S(in[5])
  );
LUT6  #(
    .INIT(64'hb7a68478e228318a)
  ) _052_ (
    .I0(in[0]),
    .I1(in[4]),
    .I2(in[3]),
    .I3(in[7]),
    .I4(in[2]),
    .I5(in[1]),
    .O(_004_)
  );
LUT6  #(
    .INIT(64'h63fa354b5e8c9feb)
  ) _053_ (
    .I0(in[0]),
    .I1(in[4]),
    .I2(in[3]),
    .I3(in[7]),
    .I4(in[2]),
    .I5(in[1]),
    .O(_005_)
  );
MUXF7  _054_ (
    .I0(_004_),
    .I1(_005_),
    .O(_001_),
    .S(in[5])
  );
MUXF8  _055_ (
    .I0(_000_),
    .I1(_001_),
    .O(_048_[0]),
    .S(in[6])
  );
LUT6  #(
    .INIT(64'h7842c7de2a355bf5)
  ) _056_ (
    .I0(in[3]),
    .I1(in[4]),
    .I2(in[2]),
    .I3(in[1]),
    .I4(in[6]),
    .I5(in[0]),
    .O(_008_)
  );
LUT6  #(
    .INIT(64'hb2587728d9abed92)
  ) _057_ (
    .I0(in[3]),
    .I1(in[4]),
    .I2(in[2]),
    .I3(in[1]),
    .I4(in[6]),
    .I5(in[0]),
    .O(_009_)
  );
MUXF7  _058_ (
    .I0(_008_),
    .I1(_009_),
    .O(_006_),
    .S(in[7])
  );
LUT6  #(
    .INIT(64'haa18f8f0195fec28)
  ) _059_ (
    .I0(in[3]),
    .I1(in[4]),
    .I2(in[2]),
    .I3(in[1]),
    .I4(in[6]),
    .I5(in[0]),
    .O(_010_)
  );
LUT6  #(
    .INIT(64'h1d612c0419bcae93)
  ) _060_ (
    .I0(in[3]),
    .I1(in[4]),
    .I2(in[2]),
    .I3(in[1]),
    .I4(in[6]),
    .I5(in[0]),
    .O(_011_)
  );
MUXF7  _061_ (
    .I0(_010_),
    .I1(_011_),
    .O(_007_),
    .S(in[7])
  );
MUXF8  _062_ (
    .I0(_006_),
    .I1(_007_),
    .O(_048_[1]),
    .S(in[5])
  );
LUT6  #(
    .INIT(64'h49d52fbbd9c93745)
  ) _063_ (
    .I0(in[3]),
    .I1(in[4]),
    .I2(in[0]),
    .I3(in[2]),
    .I4(in[5]),
    .I5(in[1]),
    .O(_014_)
  );
LUT6  #(
    .INIT(64'h8b7bc33a85d039be)
  ) _064_ (
    .I0(in[3]),
    .I1(in[4]),
    .I2(in[0]),
    .I3(in[2]),
    .I4(in[5]),
    .I5(in[1]),
    .O(_015_)
  );
MUXF7  _065_ (
    .I0(_014_),
    .I1(_015_),
    .O(_012_),
    .S(in[6])
  );
LUT6  #(
    .INIT(64'h0cb5b80790b6dda8)
  ) _066_ (
    .I0(in[3]),
    .I1(in[4]),
    .I2(in[0]),
    .I3(in[2]),
    .I4(in[5]),
    .I5(in[1]),
    .O(_016_)
  );
LUT6  #(
    .INIT(64'had82f67846225a41)
  ) _067_ (
    .I0(in[3]),
    .I1(in[4]),
    .I2(in[0]),
    .I3(in[2]),
    .I4(in[5]),
    .I5(in[1]),
    .O(_017_)
  );
MUXF7  _068_ (
    .I0(_016_),
    .I1(_017_),
    .O(_013_),
    .S(in[6])
  );
MUXF8  _069_ (
    .I0(_012_),
    .I1(_013_),
    .O(_048_[2]),
    .S(in[7])
  );
LUT6  #(
    .INIT(64'h8ff4b5ddb41a005e)
  ) _070_ (
    .I0(in[0]),
    .I1(in[4]),
    .I2(in[2]),
    .I3(in[3]),
    .I4(in[7]),
    .I5(in[1]),
    .O(_020_)
  );
LUT6  #(
    .INIT(64'h7f8b12618919a82a)
  ) _071_ (
    .I0(in[0]),
    .I1(in[4]),
    .I2(in[2]),
    .I3(in[3]),
    .I4(in[7]),
    .I5(in[1]),
    .O(_021_)
  );
MUXF7  _072_ (
    .I0(_020_),
    .I1(_021_),
    .O(_018_),
    .S(in[6])
  );
LUT6  #(
    .INIT(64'h08fceecb5f29e534)
  ) _073_ (
    .I0(in[0]),
    .I1(in[4]),
    .I2(in[2]),
    .I3(in[3]),
    .I4(in[7]),
    .I5(in[1]),
    .O(_022_)
  );
LUT6  #(
    .INIT(64'hce0de603eb2b2369)
  ) _074_ (
    .I0(in[0]),
    .I1(in[4]),
    .I2(in[2]),
    .I3(in[3]),
    .I4(in[7]),
    .I5(in[1]),
    .O(_023_)
  );
MUXF7  _075_ (
    .I0(_022_),
    .I1(_023_),
    .O(_019_),
    .S(in[6])
  );
MUXF8  _076_ (
    .I0(_018_),
    .I1(_019_),
    .O(_048_[3]),
    .S(in[5])
  );
LUT6  #(
    .INIT(64'h7fc58f6cafcd6dc4)
  ) _077_ (
    .I0(in[3]),
    .I1(in[0]),
    .I2(in[4]),
    .I3(in[6]),
    .I4(in[2]),
    .I5(in[1]),
    .O(_026_)
  );
LUT6  #(
    .INIT(64'h75321c1ab7cd444e)
  ) _078_ (
    .I0(in[3]),
    .I1(in[0]),
    .I2(in[4]),
    .I3(in[6]),
    .I4(in[2]),
    .I5(in[1]),
    .O(_027_)
  );
MUXF7  _079_ (
    .I0(_026_),
    .I1(_027_),
    .O(_024_),
    .S(in[7])
  );
LUT6  #(
    .INIT(64'hf42108eb1c54c149)
  ) _080_ (
    .I0(in[3]),
    .I1(in[0]),
    .I2(in[4]),
    .I3(in[6]),
    .I4(in[2]),
    .I5(in[1]),
    .O(_028_)
  );
LUT6  #(
    .INIT(64'h469ee26561cb493b)
  ) _081_ (
    .I0(in[3]),
    .I1(in[0]),
    .I2(in[4]),
    .I3(in[6]),
    .I4(in[2]),
    .I5(in[1]),
    .O(_029_)
  );
MUXF7  _082_ (
    .I0(_028_),
    .I1(_029_),
    .O(_025_),
    .S(in[7])
  );
MUXF8  _083_ (
    .I0(_024_),
    .I1(_025_),
    .O(_048_[4]),
    .S(in[5])
  );
LUT6  #(
    .INIT(64'hf93f687d21930b92)
  ) _084_ (
    .I0(in[0]),
    .I1(in[4]),
    .I2(in[3]),
    .I3(in[1]),
    .I4(in[5]),
    .I5(in[2]),
    .O(_032_)
  );
LUT6  #(
    .INIT(64'hddfc4d0962e5f23c)
  ) _085_ (
    .I0(in[0]),
    .I1(in[4]),
    .I2(in[3]),
    .I3(in[1]),
    .I4(in[5]),
    .I5(in[2]),
    .O(_033_)
  );
MUXF7  _086_ (
    .I0(_032_),
    .I1(_033_),
    .O(_030_),
    .S(in[6])
  );
LUT6  #(
    .INIT(64'h22b8b6e345a2f900)
  ) _087_ (
    .I0(in[0]),
    .I1(in[4]),
    .I2(in[3]),
    .I3(in[1]),
    .I4(in[5]),
    .I5(in[2]),
    .O(_034_)
  );
LUT6  #(
    .INIT(64'he2e6c52103b2f4af)
  ) _088_ (
    .I0(in[0]),
    .I1(in[4]),
    .I2(in[3]),
    .I3(in[1]),
    .I4(in[5]),
    .I5(in[2]),
    .O(_035_)
  );
MUXF7  _089_ (
    .I0(_034_),
    .I1(_035_),
    .O(_031_),
    .S(in[6])
  );
MUXF8  _090_ (
    .I0(_030_),
    .I1(_031_),
    .O(_048_[5]),
    .S(in[7])
  );
LUT6  #(
    .INIT(64'h51387b85304af57d)
  ) _091_ (
    .I0(in[4]),
    .I1(in[2]),
    .I2(in[3]),
    .I3(in[1]),
    .I4(in[7]),
    .I5(in[0]),
    .O(_038_)
  );
LUT6  #(
    .INIT(64'h2367365c1f336968)
  ) _092_ (
    .I0(in[4]),
    .I1(in[2]),
    .I2(in[3]),
    .I3(in[1]),
    .I4(in[7]),
    .I5(in[0]),
    .O(_039_)
  );
MUXF7  _093_ (
    .I0(_038_),
    .I1(_039_),
    .O(_036_),
    .S(in[6])
  );
LUT6  #(
    .INIT(64'h7a81b195f7a3d6d5)
  ) _094_ (
    .I0(in[4]),
    .I1(in[2]),
    .I2(in[3]),
    .I3(in[1]),
    .I4(in[7]),
    .I5(in[0]),
    .O(_040_)
  );
LUT6  #(
    .INIT(64'h180b79f3e08d8d20)
  ) _095_ (
    .I0(in[4]),
    .I1(in[2]),
    .I2(in[3]),
    .I3(in[1]),
    .I4(in[7]),
    .I5(in[0]),
    .O(_041_)
  );
MUXF7  _096_ (
    .I0(_040_),
    .I1(_041_),
    .O(_037_),
    .S(in[6])
  );
MUXF8  _097_ (
    .I0(_036_),
    .I1(_037_),
    .O(_048_[6]),
    .S(in[5])
  );
LUT6  #(
    .INIT(64'h89ab56b3fd5f5795)
  ) _098_ (
    .I0(in[3]),
    .I1(in[0]),
    .I2(in[4]),
    .I3(in[1]),
    .I4(in[2]),
    .I5(in[7]),
    .O(_044_)
  );
LUT6  #(
    .INIT(64'h1ee1e8fb852aca44)
  ) _099_ (
    .I0(in[3]),
    .I1(in[0]),
    .I2(in[4]),
    .I3(in[1]),
    .I4(in[2]),
    .I5(in[7]),
    .O(_045_)
  );
MUXF7  _100_ (
    .I0(_044_),
    .I1(_045_),
    .O(_042_),
    .S(in[5])
  );
LUT6  #(
    .INIT(64'h1492623ee1ec42f2)
  ) _101_ (
    .I0(in[3]),
    .I1(in[0]),
    .I2(in[4]),
    .I3(in[1]),
    .I4(in[2]),
    .I5(in[7]),
    .O(_046_)
  );
LUT6  #(
    .INIT(64'h58cf0825e0873c1f)
  ) _102_ (
    .I0(in[3]),
    .I1(in[0]),
    .I2(in[4]),
    .I3(in[1]),
    .I4(in[2]),
    .I5(in[7]),
    .O(_047_)
  );
MUXF7  _103_ (
    .I0(_046_),
    .I1(_047_),
    .O(_043_),
    .S(in[5])
  );
MUXF8  _104_ (
    .I0(_042_),
    .I1(_043_),
    .O(_048_[7]),
    .S(in[6])
  );
FDRE  #(
    .INIT(1'hx)
  ) _105_ (
    .C(clk),
    .CE(1'h1),
    .D(_048_[0]),
    .Q(out[0]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _106_ (
    .C(clk),
    .CE(1'h1),
    .D(_048_[1]),
    .Q(out[1]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _107_ (
    .C(clk),
    .CE(1'h1),
    .D(_048_[2]),
    .Q(out[2]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _108_ (
    .C(clk),
    .CE(1'h1),
    .D(_048_[3]),
    .Q(out[3]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _109_ (
    .C(clk),
    .CE(1'h1),
    .D(_048_[4]),
    .Q(out[4]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _110_ (
    .C(clk),
    .CE(1'h1),
    .D(_048_[5]),
    .Q(out[5]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _111_ (
    .C(clk),
    .CE(1'h1),
    .D(_048_[6]),
    .Q(out[6]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _112_ (
    .C(clk),
    .CE(1'h1),
    .D(_048_[7]),
    .Q(out[7]),
    .R(1'h0)
  );
endmodule
