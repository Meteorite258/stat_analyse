module wb_conmax_top(clk_i,  rst_i, m0_data_i, m0_data_o, m0_addr_i, m0_sel_i, m0_we_i, m0_cyc_i, m0_stb_i, m0_ack_o, m0_err_o, m0_rty_o, m1_data_i, m1_data_o, m1_addr_i, m1_sel_i, m1_we_i, m1_cyc_i, m1_stb_i, m1_ack_o, m1_err_o
, m1_rty_o, m2_data_i, m2_data_o, m2_addr_i, m2_sel_i, m2_we_i, m2_cyc_i, m2_stb_i, m2_ack_o, m2_err_o, m2_rty_o, m3_data_i, m3_data_o, m3_addr_i, m3_sel_i, m3_we_i, m3_cyc_i, m3_stb_i, m3_ack_o, m3_err_o, m3_rty_o
, m4_data_i, m4_data_o, m4_addr_i, m4_sel_i, m4_we_i, m4_cyc_i, m4_stb_i, m4_ack_o, m4_err_o, m4_rty_o, m5_data_i, m5_data_o, m5_addr_i, m5_sel_i, m5_we_i, m5_cyc_i, m5_stb_i, m5_ack_o, m5_err_o, m5_rty_o, m6_data_i
, m6_data_o, m6_addr_i, m6_sel_i, m6_we_i, m6_cyc_i, m6_stb_i, m6_ack_o, m6_err_o, m6_rty_o, m7_data_i, m7_data_o, m7_addr_i, m7_sel_i, m7_we_i, m7_cyc_i, m7_stb_i, m7_ack_o, m7_err_o, m7_rty_o, s0_data_i, s0_data_o
, s0_addr_o, s0_sel_o, s0_we_o, s0_cyc_o, s0_stb_o, s0_ack_i, s0_err_i, s0_rty_i, s1_data_i, s1_data_o, s1_addr_o, s1_sel_o, s1_we_o, s1_cyc_o, s1_stb_o, s1_ack_i, s1_err_i, s1_rty_i, s2_data_i, s2_data_o, s2_addr_o
, s2_sel_o, s2_we_o, s2_cyc_o, s2_stb_o, s2_ack_i, s2_err_i, s2_rty_i, s3_data_i, s3_data_o, s3_addr_o, s3_sel_o, s3_we_o, s3_cyc_o, s3_stb_o, s3_ack_i, s3_err_i, s3_rty_i, s4_data_i, s4_data_o, s4_addr_o, s4_sel_o
, s4_we_o, s4_cyc_o, s4_stb_o, s4_ack_i, s4_err_i, s4_rty_i, s5_data_i, s5_data_o, s5_addr_o, s5_sel_o, s5_we_o, s5_cyc_o, s5_stb_o, s5_ack_i, s5_err_i, s5_rty_i, s6_data_i, s6_data_o, s6_addr_o, s6_sel_o, s6_we_o
, s6_cyc_o, s6_stb_o, s6_ack_i, s6_err_i, s6_rty_i, s7_data_i, s7_data_o, s7_addr_o, s7_sel_o, s7_we_o, s7_cyc_o, s7_stb_o, s7_ack_i, s7_err_i, s7_rty_i, s8_data_i, s8_data_o, s8_addr_o, s8_sel_o, s8_we_o, s8_cyc_o
, s8_stb_o, s8_ack_i, s8_err_i, s8_rty_i, s9_data_i, s9_data_o, s9_addr_o, s9_sel_o, s9_we_o, s9_cyc_o, s9_stb_o, s9_ack_i, s9_err_i, s9_rty_i, s10_data_i, s10_data_o, s10_addr_o, s10_sel_o, s10_we_o, s10_cyc_o, s10_stb_o
, s10_ack_i, s10_err_i, s10_rty_i, s11_data_i, s11_data_o, s11_addr_o, s11_sel_o, s11_we_o, s11_cyc_o, s11_stb_o, s11_ack_i, s11_err_i, s11_rty_i, s12_data_i, s12_data_o, s12_addr_o, s12_sel_o, s12_we_o, s12_cyc_o, s12_stb_o, s12_ack_i
, s12_err_i, s12_rty_i, s13_data_i, s13_data_o, s13_addr_o, s13_sel_o, s13_we_o, s13_cyc_o, s13_stb_o, s13_ack_i, s13_err_i, s13_rty_i, s14_data_i, s14_data_o, s14_addr_o, s14_sel_o, s14_we_o, s14_cyc_o, s14_stb_o, s14_ack_i, s14_err_i
, s14_rty_i, s15_data_i, s15_data_o, s15_addr_o, s15_sel_o, s15_we_o, s15_cyc_o, s15_stb_o, s15_ack_i, s15_err_i, s15_rty_i);
wire  _0000_;
wire  _0001_;
wire  _0002_;
wire  [31:0] _0003_;
wire  _0004_;
wire  [31:0] _0005_;
wire  [31:0] _0006_;
wire  _0007_;
wire  _0008_;
wire  [3:0] _0009_;
wire  _0010_;
wire  _0011_;
wire  _0012_;
wire  [31:0] _0013_;
wire  _0014_;
wire  [31:0] _0015_;
wire  [31:0] _0016_;
wire  _0017_;
wire  _0018_;
wire  [3:0] _0019_;
wire  _0020_;
wire  _0021_;
wire  _0022_;
wire  [31:0] _0023_;
wire  _0024_;
wire  [31:0] _0025_;
wire  [31:0] _0026_;
wire  _0027_;
wire  _0028_;
wire  [3:0] _0029_;
wire  _0030_;
wire  _0031_;
wire  _0032_;
wire  [31:0] _0033_;
wire  _0034_;
wire  [31:0] _0035_;
wire  [31:0] _0036_;
wire  _0037_;
wire  _0038_;
wire  [3:0] _0039_;
wire  _0040_;
wire  _0041_;
wire  _0042_;
wire  [31:0] _0043_;
wire  _0044_;
wire  [31:0] _0045_;
wire  [31:0] _0046_;
wire  _0047_;
wire  _0048_;
wire  [3:0] _0049_;
wire  _0050_;
wire  _0051_;
wire  _0052_;
wire  [31:0] _0053_;
wire  _0054_;
wire  [31:0] _0055_;
wire  [31:0] _0056_;
wire  _0057_;
wire  _0058_;
wire  [3:0] _0059_;
wire  _0060_;
wire  _0061_;
wire  _0062_;
wire  [31:0] _0063_;
wire  _0064_;
wire  [31:0] _0065_;
wire  [31:0] _0066_;
wire  _0067_;
wire  _0068_;
wire  [3:0] _0069_;
wire  _0070_;
wire  _0071_;
wire  _0072_;
wire  [31:0] _0073_;
wire  _0074_;
wire  [31:0] _0075_;
wire  [31:0] _0076_;
wire  _0077_;
wire  _0078_;
wire  [3:0] _0079_;
wire  _0080_;
wire  _0081_;
wire  _0082_;
wire  _0083_;
wire  [31:0] _0084_;
wire  _0085_;
wire  [31:0] _0086_;
wire  [31:0] _0087_;
wire  _0088_;
wire  _0089_;
wire  [3:0] _0090_;
wire  _0091_;
wire  _0092_;
wire  _0093_;
wire  [31:0] _0094_;
wire  _0095_;
wire  [31:0] _0096_;
wire  [31:0] _0097_;
wire  _0098_;
wire  _0099_;
wire  [3:0] _0100_;
wire  _0101_;
wire  _0102_;
wire  _0103_;
wire  [31:0] _0104_;
wire  _0105_;
wire  [31:0] _0106_;
wire  [31:0] _0107_;
wire  _0108_;
wire  _0109_;
wire  [3:0] _0110_;
wire  _0111_;
wire  _0112_;
wire  _0113_;
wire  [31:0] _0114_;
wire  _0115_;
wire  [31:0] _0116_;
wire  [31:0] _0117_;
wire  _0118_;
wire  _0119_;
wire  [3:0] _0120_;
wire  _0121_;
wire  _0122_;
wire  _0123_;
wire  [31:0] _0124_;
wire  _0125_;
wire  [31:0] _0126_;
wire  [31:0] _0127_;
wire  _0128_;
wire  _0129_;
wire  [3:0] _0130_;
wire  _0131_;
wire  _0132_;
wire  _0133_;
wire  [31:0] _0134_;
wire  _0135_;
wire  [31:0] _0136_;
wire  [31:0] _0137_;
wire  _0138_;
wire  _0139_;
wire  [3:0] _0140_;
wire  _0141_;
wire  _0142_;
wire  _0143_;
wire  [31:0] _0144_;
wire  _0145_;
wire  [31:0] _0146_;
wire  [31:0] _0147_;
wire  _0148_;
wire  _0149_;
wire  [3:0] _0150_;
wire  _0151_;
wire  _0152_;
wire  _0153_;
wire  [31:0] _0154_;
wire  _0155_;
wire  [31:0] _0156_;
wire  [31:0] _0157_;
wire  _0158_;
wire  _0159_;
wire  [3:0] _0160_;
wire  _0161_;
wire  _0162_;
wire  _0163_;
wire  [31:0] _0164_;
wire  _0165_;
wire  [31:0] _0166_;
wire  [31:0] _0167_;
wire  _0168_;
wire  _0169_;
wire  [3:0] _0170_;
wire  _0171_;
wire  _0172_;
wire  _0173_;
wire  [31:0] _0174_;
wire  _0175_;
wire  [31:0] _0176_;
wire  [31:0] _0177_;
wire  _0178_;
wire  _0179_;
wire  [3:0] _0180_;
wire  _0181_;
wire  _0182_;
wire  _0183_;
wire  [31:0] _0184_;
wire  _0185_;
wire  [31:0] _0186_;
wire  [31:0] _0187_;
wire  _0188_;
wire  _0189_;
wire  [3:0] _0190_;
wire  _0191_;
wire  _0192_;
wire  _0193_;
wire  [31:0] _0194_;
wire  _0195_;
wire  [31:0] _0196_;
wire  [31:0] _0197_;
wire  _0198_;
wire  _0199_;
wire  [3:0] _0200_;
wire  _0201_;
wire  _0202_;
wire  _0203_;
wire  [31:0] _0204_;
wire  _0205_;
wire  [31:0] _0206_;
wire  [31:0] _0207_;
wire  _0208_;
wire  _0209_;
wire  [3:0] _0210_;
wire  _0211_;
wire  _0212_;
wire  _0213_;
wire  [31:0] _0214_;
wire  _0215_;
wire  [31:0] _0216_;
wire  [31:0] _0217_;
wire  _0218_;
wire  _0219_;
wire  [3:0] _0220_;
wire  _0221_;
wire  _0222_;
wire  _0223_;
wire  [31:0] _0224_;
wire  _0225_;
wire  [31:0] _0226_;
wire  [31:0] _0227_;
wire  _0228_;
wire  _0229_;
wire  [3:0] _0230_;
wire  _0231_;
wire  _0232_;
wire  _0233_;
wire  [31:0] _0234_;
wire  _0235_;
wire  [31:0] _0236_;
wire  [31:0] _0237_;
wire  _0238_;
wire  _0239_;
wire  [3:0] _0240_;
wire  _0241_;
wire  _0242_;
input  clk_i;
wire  clk_i;
wire  [15:0] conf0;
wire  [15:0] conf1;
wire  [15:0] conf10;
wire  [15:0] conf11;
wire  [15:0] conf12;
wire  [15:0] conf13;
wire  [15:0] conf14;
wire  [15:0] conf15;
wire  [15:0] conf2;
wire  [15:0] conf3;
wire  [15:0] conf4;
wire  [15:0] conf5;
wire  [15:0] conf6;
wire  [15:0] conf7;
wire  [15:0] conf8;
wire  [15:0] conf9;
wire  i_s15_ack_i;
wire  [31:0] i_s15_addr_o;
wire  i_s15_cyc_o;
wire  [31:0] i_s15_data_i;
wire  [31:0] i_s15_data_o;
wire  i_s15_err_i;
wire  i_s15_rty_i;
wire  [3:0] i_s15_sel_o;
wire  i_s15_stb_o;
wire  i_s15_we_o;
output  m0_ack_o;
wire  m0_ack_o;
input  [31:0] m0_addr_i;
wire  [31:0] m0_addr_i;
input  m0_cyc_i;
wire  m0_cyc_i;
input  [31:0] m0_data_i;
wire  [31:0] m0_data_i;
output  [31:0] m0_data_o;
wire  [31:0] m0_data_o;
output  m0_err_o;
wire  m0_err_o;
output  m0_rty_o;
wire  m0_rty_o;
input  [3:0] m0_sel_i;
wire  [3:0] m0_sel_i;
input  m0_stb_i;
wire  m0_stb_i;
input  m0_we_i;
wire  m0_we_i;
wire  m0s0_ack;
wire  [31:0] m0s0_addr;
wire  m0s0_cyc;
wire  [31:0] m0s0_data_i;
wire  [31:0] m0s0_data_o;
wire  m0s0_err;
wire  m0s0_rty;
wire  [3:0] m0s0_sel;
wire  m0s0_stb;
wire  m0s0_we;
wire  m0s10_ack;
wire  [31:0] m0s10_addr;
wire  m0s10_cyc;
wire  [31:0] m0s10_data_i;
wire  [31:0] m0s10_data_o;
wire  m0s10_err;
wire  m0s10_rty;
wire  [3:0] m0s10_sel;
wire  m0s10_stb;
wire  m0s10_we;
wire  m0s11_ack;
wire  [31:0] m0s11_addr;
wire  m0s11_cyc;
wire  [31:0] m0s11_data_i;
wire  [31:0] m0s11_data_o;
wire  m0s11_err;
wire  m0s11_rty;
wire  [3:0] m0s11_sel;
wire  m0s11_stb;
wire  m0s11_we;
wire  m0s12_ack;
wire  [31:0] m0s12_addr;
wire  m0s12_cyc;
wire  [31:0] m0s12_data_i;
wire  [31:0] m0s12_data_o;
wire  m0s12_err;
wire  m0s12_rty;
wire  [3:0] m0s12_sel;
wire  m0s12_stb;
wire  m0s12_we;
wire  m0s13_ack;
wire  [31:0] m0s13_addr;
wire  m0s13_cyc;
wire  [31:0] m0s13_data_i;
wire  [31:0] m0s13_data_o;
wire  m0s13_err;
wire  m0s13_rty;
wire  [3:0] m0s13_sel;
wire  m0s13_stb;
wire  m0s13_we;
wire  m0s14_ack;
wire  [31:0] m0s14_addr;
wire  m0s14_cyc;
wire  [31:0] m0s14_data_i;
wire  [31:0] m0s14_data_o;
wire  m0s14_err;
wire  m0s14_rty;
wire  [3:0] m0s14_sel;
wire  m0s14_stb;
wire  m0s14_we;
wire  m0s15_ack;
wire  [31:0] m0s15_addr;
wire  m0s15_cyc;
wire  [31:0] m0s15_data_i;
wire  [31:0] m0s15_data_o;
wire  m0s15_err;
wire  m0s15_rty;
wire  [3:0] m0s15_sel;
wire  m0s15_stb;
wire  m0s15_we;
wire  m0s1_ack;
wire  [31:0] m0s1_addr;
wire  m0s1_cyc;
wire  [31:0] m0s1_data_i;
wire  [31:0] m0s1_data_o;
wire  m0s1_err;
wire  m0s1_rty;
wire  [3:0] m0s1_sel;
wire  m0s1_stb;
wire  m0s1_we;
wire  m0s2_ack;
wire  [31:0] m0s2_addr;
wire  m0s2_cyc;
wire  [31:0] m0s2_data_i;
wire  [31:0] m0s2_data_o;
wire  m0s2_err;
wire  m0s2_rty;
wire  [3:0] m0s2_sel;
wire  m0s2_stb;
wire  m0s2_we;
wire  m0s3_ack;
wire  [31:0] m0s3_addr;
wire  m0s3_cyc;
wire  [31:0] m0s3_data_i;
wire  [31:0] m0s3_data_o;
wire  m0s3_err;
wire  m0s3_rty;
wire  [3:0] m0s3_sel;
wire  m0s3_stb;
wire  m0s3_we;
wire  m0s4_ack;
wire  [31:0] m0s4_addr;
wire  m0s4_cyc;
wire  [31:0] m0s4_data_i;
wire  [31:0] m0s4_data_o;
wire  m0s4_err;
wire  m0s4_rty;
wire  [3:0] m0s4_sel;
wire  m0s4_stb;
wire  m0s4_we;
wire  m0s5_ack;
wire  [31:0] m0s5_addr;
wire  m0s5_cyc;
wire  [31:0] m0s5_data_i;
wire  [31:0] m0s5_data_o;
wire  m0s5_err;
wire  m0s5_rty;
wire  [3:0] m0s5_sel;
wire  m0s5_stb;
wire  m0s5_we;
wire  m0s6_ack;
wire  [31:0] m0s6_addr;
wire  m0s6_cyc;
wire  [31:0] m0s6_data_i;
wire  [31:0] m0s6_data_o;
wire  m0s6_err;
wire  m0s6_rty;
wire  [3:0] m0s6_sel;
wire  m0s6_stb;
wire  m0s6_we;
wire  m0s7_ack;
wire  [31:0] m0s7_addr;
wire  m0s7_cyc;
wire  [31:0] m0s7_data_i;
wire  [31:0] m0s7_data_o;
wire  m0s7_err;
wire  m0s7_rty;
wire  [3:0] m0s7_sel;
wire  m0s7_stb;
wire  m0s7_we;
wire  m0s8_ack;
wire  [31:0] m0s8_addr;
wire  m0s8_cyc;
wire  [31:0] m0s8_data_i;
wire  [31:0] m0s8_data_o;
wire  m0s8_err;
wire  m0s8_rty;
wire  [3:0] m0s8_sel;
wire  m0s8_stb;
wire  m0s8_we;
wire  m0s9_ack;
wire  [31:0] m0s9_addr;
wire  m0s9_cyc;
wire  [31:0] m0s9_data_i;
wire  [31:0] m0s9_data_o;
wire  m0s9_err;
wire  m0s9_rty;
wire  [3:0] m0s9_sel;
wire  m0s9_stb;
wire  m0s9_we;
output  m1_ack_o;
wire  m1_ack_o;
input  [31:0] m1_addr_i;
wire  [31:0] m1_addr_i;
input  m1_cyc_i;
wire  m1_cyc_i;
input  [31:0] m1_data_i;
wire  [31:0] m1_data_i;
output  [31:0] m1_data_o;
wire  [31:0] m1_data_o;
output  m1_err_o;
wire  m1_err_o;
output  m1_rty_o;
wire  m1_rty_o;
input  [3:0] m1_sel_i;
wire  [3:0] m1_sel_i;
input  m1_stb_i;
wire  m1_stb_i;
input  m1_we_i;
wire  m1_we_i;
wire  m1s0_ack;
wire  [31:0] m1s0_addr;
wire  m1s0_cyc;
wire  [31:0] m1s0_data_i;
wire  [31:0] m1s0_data_o;
wire  m1s0_err;
wire  m1s0_rty;
wire  [3:0] m1s0_sel;
wire  m1s0_stb;
wire  m1s0_we;
wire  m1s10_ack;
wire  [31:0] m1s10_addr;
wire  m1s10_cyc;
wire  [31:0] m1s10_data_i;
wire  [31:0] m1s10_data_o;
wire  m1s10_err;
wire  m1s10_rty;
wire  [3:0] m1s10_sel;
wire  m1s10_stb;
wire  m1s10_we;
wire  m1s11_ack;
wire  [31:0] m1s11_addr;
wire  m1s11_cyc;
wire  [31:0] m1s11_data_i;
wire  [31:0] m1s11_data_o;
wire  m1s11_err;
wire  m1s11_rty;
wire  [3:0] m1s11_sel;
wire  m1s11_stb;
wire  m1s11_we;
wire  m1s12_ack;
wire  [31:0] m1s12_addr;
wire  m1s12_cyc;
wire  [31:0] m1s12_data_i;
wire  [31:0] m1s12_data_o;
wire  m1s12_err;
wire  m1s12_rty;
wire  [3:0] m1s12_sel;
wire  m1s12_stb;
wire  m1s12_we;
wire  m1s13_ack;
wire  [31:0] m1s13_addr;
wire  m1s13_cyc;
wire  [31:0] m1s13_data_i;
wire  [31:0] m1s13_data_o;
wire  m1s13_err;
wire  m1s13_rty;
wire  [3:0] m1s13_sel;
wire  m1s13_stb;
wire  m1s13_we;
wire  m1s14_ack;
wire  [31:0] m1s14_addr;
wire  m1s14_cyc;
wire  [31:0] m1s14_data_i;
wire  [31:0] m1s14_data_o;
wire  m1s14_err;
wire  m1s14_rty;
wire  [3:0] m1s14_sel;
wire  m1s14_stb;
wire  m1s14_we;
wire  m1s15_ack;
wire  [31:0] m1s15_addr;
wire  m1s15_cyc;
wire  [31:0] m1s15_data_i;
wire  [31:0] m1s15_data_o;
wire  m1s15_err;
wire  m1s15_rty;
wire  [3:0] m1s15_sel;
wire  m1s15_stb;
wire  m1s15_we;
wire  m1s1_ack;
wire  [31:0] m1s1_addr;
wire  m1s1_cyc;
wire  [31:0] m1s1_data_i;
wire  [31:0] m1s1_data_o;
wire  m1s1_err;
wire  m1s1_rty;
wire  [3:0] m1s1_sel;
wire  m1s1_stb;
wire  m1s1_we;
wire  m1s2_ack;
wire  [31:0] m1s2_addr;
wire  m1s2_cyc;
wire  [31:0] m1s2_data_i;
wire  [31:0] m1s2_data_o;
wire  m1s2_err;
wire  m1s2_rty;
wire  [3:0] m1s2_sel;
wire  m1s2_stb;
wire  m1s2_we;
wire  m1s3_ack;
wire  [31:0] m1s3_addr;
wire  m1s3_cyc;
wire  [31:0] m1s3_data_i;
wire  [31:0] m1s3_data_o;
wire  m1s3_err;
wire  m1s3_rty;
wire  [3:0] m1s3_sel;
wire  m1s3_stb;
wire  m1s3_we;
wire  m1s4_ack;
wire  [31:0] m1s4_addr;
wire  m1s4_cyc;
wire  [31:0] m1s4_data_i;
wire  [31:0] m1s4_data_o;
wire  m1s4_err;
wire  m1s4_rty;
wire  [3:0] m1s4_sel;
wire  m1s4_stb;
wire  m1s4_we;
wire  m1s5_ack;
wire  [31:0] m1s5_addr;
wire  m1s5_cyc;
wire  [31:0] m1s5_data_i;
wire  [31:0] m1s5_data_o;
wire  m1s5_err;
wire  m1s5_rty;
wire  [3:0] m1s5_sel;
wire  m1s5_stb;
wire  m1s5_we;
wire  m1s6_ack;
wire  [31:0] m1s6_addr;
wire  m1s6_cyc;
wire  [31:0] m1s6_data_i;
wire  [31:0] m1s6_data_o;
wire  m1s6_err;
wire  m1s6_rty;
wire  [3:0] m1s6_sel;
wire  m1s6_stb;
wire  m1s6_we;
wire  m1s7_ack;
wire  [31:0] m1s7_addr;
wire  m1s7_cyc;
wire  [31:0] m1s7_data_i;
wire  [31:0] m1s7_data_o;
wire  m1s7_err;
wire  m1s7_rty;
wire  [3:0] m1s7_sel;
wire  m1s7_stb;
wire  m1s7_we;
wire  m1s8_ack;
wire  [31:0] m1s8_addr;
wire  m1s8_cyc;
wire  [31:0] m1s8_data_i;
wire  [31:0] m1s8_data_o;
wire  m1s8_err;
wire  m1s8_rty;
wire  [3:0] m1s8_sel;
wire  m1s8_stb;
wire  m1s8_we;
wire  m1s9_ack;
wire  [31:0] m1s9_addr;
wire  m1s9_cyc;
wire  [31:0] m1s9_data_i;
wire  [31:0] m1s9_data_o;
wire  m1s9_err;
wire  m1s9_rty;
wire  [3:0] m1s9_sel;
wire  m1s9_stb;
wire  m1s9_we;
output  m2_ack_o;
wire  m2_ack_o;
input  [31:0] m2_addr_i;
wire  [31:0] m2_addr_i;
input  m2_cyc_i;
wire  m2_cyc_i;
input  [31:0] m2_data_i;
wire  [31:0] m2_data_i;
output  [31:0] m2_data_o;
wire  [31:0] m2_data_o;
output  m2_err_o;
wire  m2_err_o;
output  m2_rty_o;
wire  m2_rty_o;
input  [3:0] m2_sel_i;
wire  [3:0] m2_sel_i;
input  m2_stb_i;
wire  m2_stb_i;
input  m2_we_i;
wire  m2_we_i;
wire  m2s0_ack;
wire  [31:0] m2s0_addr;
wire  m2s0_cyc;
wire  [31:0] m2s0_data_i;
wire  [31:0] m2s0_data_o;
wire  m2s0_err;
wire  m2s0_rty;
wire  [3:0] m2s0_sel;
wire  m2s0_stb;
wire  m2s0_we;
wire  m2s10_ack;
wire  [31:0] m2s10_addr;
wire  m2s10_cyc;
wire  [31:0] m2s10_data_i;
wire  [31:0] m2s10_data_o;
wire  m2s10_err;
wire  m2s10_rty;
wire  [3:0] m2s10_sel;
wire  m2s10_stb;
wire  m2s10_we;
wire  m2s11_ack;
wire  [31:0] m2s11_addr;
wire  m2s11_cyc;
wire  [31:0] m2s11_data_i;
wire  [31:0] m2s11_data_o;
wire  m2s11_err;
wire  m2s11_rty;
wire  [3:0] m2s11_sel;
wire  m2s11_stb;
wire  m2s11_we;
wire  m2s12_ack;
wire  [31:0] m2s12_addr;
wire  m2s12_cyc;
wire  [31:0] m2s12_data_i;
wire  [31:0] m2s12_data_o;
wire  m2s12_err;
wire  m2s12_rty;
wire  [3:0] m2s12_sel;
wire  m2s12_stb;
wire  m2s12_we;
wire  m2s13_ack;
wire  [31:0] m2s13_addr;
wire  m2s13_cyc;
wire  [31:0] m2s13_data_i;
wire  [31:0] m2s13_data_o;
wire  m2s13_err;
wire  m2s13_rty;
wire  [3:0] m2s13_sel;
wire  m2s13_stb;
wire  m2s13_we;
wire  m2s14_ack;
wire  [31:0] m2s14_addr;
wire  m2s14_cyc;
wire  [31:0] m2s14_data_i;
wire  [31:0] m2s14_data_o;
wire  m2s14_err;
wire  m2s14_rty;
wire  [3:0] m2s14_sel;
wire  m2s14_stb;
wire  m2s14_we;
wire  m2s15_ack;
wire  [31:0] m2s15_addr;
wire  m2s15_cyc;
wire  [31:0] m2s15_data_i;
wire  [31:0] m2s15_data_o;
wire  m2s15_err;
wire  m2s15_rty;
wire  [3:0] m2s15_sel;
wire  m2s15_stb;
wire  m2s15_we;
wire  m2s1_ack;
wire  [31:0] m2s1_addr;
wire  m2s1_cyc;
wire  [31:0] m2s1_data_i;
wire  [31:0] m2s1_data_o;
wire  m2s1_err;
wire  m2s1_rty;
wire  [3:0] m2s1_sel;
wire  m2s1_stb;
wire  m2s1_we;
wire  m2s2_ack;
wire  [31:0] m2s2_addr;
wire  m2s2_cyc;
wire  [31:0] m2s2_data_i;
wire  [31:0] m2s2_data_o;
wire  m2s2_err;
wire  m2s2_rty;
wire  [3:0] m2s2_sel;
wire  m2s2_stb;
wire  m2s2_we;
wire  m2s3_ack;
wire  [31:0] m2s3_addr;
wire  m2s3_cyc;
wire  [31:0] m2s3_data_i;
wire  [31:0] m2s3_data_o;
wire  m2s3_err;
wire  m2s3_rty;
wire  [3:0] m2s3_sel;
wire  m2s3_stb;
wire  m2s3_we;
wire  m2s4_ack;
wire  [31:0] m2s4_addr;
wire  m2s4_cyc;
wire  [31:0] m2s4_data_i;
wire  [31:0] m2s4_data_o;
wire  m2s4_err;
wire  m2s4_rty;
wire  [3:0] m2s4_sel;
wire  m2s4_stb;
wire  m2s4_we;
wire  m2s5_ack;
wire  [31:0] m2s5_addr;
wire  m2s5_cyc;
wire  [31:0] m2s5_data_i;
wire  [31:0] m2s5_data_o;
wire  m2s5_err;
wire  m2s5_rty;
wire  [3:0] m2s5_sel;
wire  m2s5_stb;
wire  m2s5_we;
wire  m2s6_ack;
wire  [31:0] m2s6_addr;
wire  m2s6_cyc;
wire  [31:0] m2s6_data_i;
wire  [31:0] m2s6_data_o;
wire  m2s6_err;
wire  m2s6_rty;
wire  [3:0] m2s6_sel;
wire  m2s6_stb;
wire  m2s6_we;
wire  m2s7_ack;
wire  [31:0] m2s7_addr;
wire  m2s7_cyc;
wire  [31:0] m2s7_data_i;
wire  [31:0] m2s7_data_o;
wire  m2s7_err;
wire  m2s7_rty;
wire  [3:0] m2s7_sel;
wire  m2s7_stb;
wire  m2s7_we;
wire  m2s8_ack;
wire  [31:0] m2s8_addr;
wire  m2s8_cyc;
wire  [31:0] m2s8_data_i;
wire  [31:0] m2s8_data_o;
wire  m2s8_err;
wire  m2s8_rty;
wire  [3:0] m2s8_sel;
wire  m2s8_stb;
wire  m2s8_we;
wire  m2s9_ack;
wire  [31:0] m2s9_addr;
wire  m2s9_cyc;
wire  [31:0] m2s9_data_i;
wire  [31:0] m2s9_data_o;
wire  m2s9_err;
wire  m2s9_rty;
wire  [3:0] m2s9_sel;
wire  m2s9_stb;
wire  m2s9_we;
output  m3_ack_o;
wire  m3_ack_o;
input  [31:0] m3_addr_i;
wire  [31:0] m3_addr_i;
input  m3_cyc_i;
wire  m3_cyc_i;
input  [31:0] m3_data_i;
wire  [31:0] m3_data_i;
output  [31:0] m3_data_o;
wire  [31:0] m3_data_o;
output  m3_err_o;
wire  m3_err_o;
output  m3_rty_o;
wire  m3_rty_o;
input  [3:0] m3_sel_i;
wire  [3:0] m3_sel_i;
input  m3_stb_i;
wire  m3_stb_i;
input  m3_we_i;
wire  m3_we_i;
wire  m3s0_ack;
wire  [31:0] m3s0_addr;
wire  m3s0_cyc;
wire  [31:0] m3s0_data_i;
wire  [31:0] m3s0_data_o;
wire  m3s0_err;
wire  m3s0_rty;
wire  [3:0] m3s0_sel;
wire  m3s0_stb;
wire  m3s0_we;
wire  m3s10_ack;
wire  [31:0] m3s10_addr;
wire  m3s10_cyc;
wire  [31:0] m3s10_data_i;
wire  [31:0] m3s10_data_o;
wire  m3s10_err;
wire  m3s10_rty;
wire  [3:0] m3s10_sel;
wire  m3s10_stb;
wire  m3s10_we;
wire  m3s11_ack;
wire  [31:0] m3s11_addr;
wire  m3s11_cyc;
wire  [31:0] m3s11_data_i;
wire  [31:0] m3s11_data_o;
wire  m3s11_err;
wire  m3s11_rty;
wire  [3:0] m3s11_sel;
wire  m3s11_stb;
wire  m3s11_we;
wire  m3s12_ack;
wire  [31:0] m3s12_addr;
wire  m3s12_cyc;
wire  [31:0] m3s12_data_i;
wire  [31:0] m3s12_data_o;
wire  m3s12_err;
wire  m3s12_rty;
wire  [3:0] m3s12_sel;
wire  m3s12_stb;
wire  m3s12_we;
wire  m3s13_ack;
wire  [31:0] m3s13_addr;
wire  m3s13_cyc;
wire  [31:0] m3s13_data_i;
wire  [31:0] m3s13_data_o;
wire  m3s13_err;
wire  m3s13_rty;
wire  [3:0] m3s13_sel;
wire  m3s13_stb;
wire  m3s13_we;
wire  m3s14_ack;
wire  [31:0] m3s14_addr;
wire  m3s14_cyc;
wire  [31:0] m3s14_data_i;
wire  [31:0] m3s14_data_o;
wire  m3s14_err;
wire  m3s14_rty;
wire  [3:0] m3s14_sel;
wire  m3s14_stb;
wire  m3s14_we;
wire  m3s15_ack;
wire  [31:0] m3s15_addr;
wire  m3s15_cyc;
wire  [31:0] m3s15_data_i;
wire  [31:0] m3s15_data_o;
wire  m3s15_err;
wire  m3s15_rty;
wire  [3:0] m3s15_sel;
wire  m3s15_stb;
wire  m3s15_we;
wire  m3s1_ack;
wire  [31:0] m3s1_addr;
wire  m3s1_cyc;
wire  [31:0] m3s1_data_i;
wire  [31:0] m3s1_data_o;
wire  m3s1_err;
wire  m3s1_rty;
wire  [3:0] m3s1_sel;
wire  m3s1_stb;
wire  m3s1_we;
wire  m3s2_ack;
wire  [31:0] m3s2_addr;
wire  m3s2_cyc;
wire  [31:0] m3s2_data_i;
wire  [31:0] m3s2_data_o;
wire  m3s2_err;
wire  m3s2_rty;
wire  [3:0] m3s2_sel;
wire  m3s2_stb;
wire  m3s2_we;
wire  m3s3_ack;
wire  [31:0] m3s3_addr;
wire  m3s3_cyc;
wire  [31:0] m3s3_data_i;
wire  [31:0] m3s3_data_o;
wire  m3s3_err;
wire  m3s3_rty;
wire  [3:0] m3s3_sel;
wire  m3s3_stb;
wire  m3s3_we;
wire  m3s4_ack;
wire  [31:0] m3s4_addr;
wire  m3s4_cyc;
wire  [31:0] m3s4_data_i;
wire  [31:0] m3s4_data_o;
wire  m3s4_err;
wire  m3s4_rty;
wire  [3:0] m3s4_sel;
wire  m3s4_stb;
wire  m3s4_we;
wire  m3s5_ack;
wire  [31:0] m3s5_addr;
wire  m3s5_cyc;
wire  [31:0] m3s5_data_i;
wire  [31:0] m3s5_data_o;
wire  m3s5_err;
wire  m3s5_rty;
wire  [3:0] m3s5_sel;
wire  m3s5_stb;
wire  m3s5_we;
wire  m3s6_ack;
wire  [31:0] m3s6_addr;
wire  m3s6_cyc;
wire  [31:0] m3s6_data_i;
wire  [31:0] m3s6_data_o;
wire  m3s6_err;
wire  m3s6_rty;
wire  [3:0] m3s6_sel;
wire  m3s6_stb;
wire  m3s6_we;
wire  m3s7_ack;
wire  [31:0] m3s7_addr;
wire  m3s7_cyc;
wire  [31:0] m3s7_data_i;
wire  [31:0] m3s7_data_o;
wire  m3s7_err;
wire  m3s7_rty;
wire  [3:0] m3s7_sel;
wire  m3s7_stb;
wire  m3s7_we;
wire  m3s8_ack;
wire  [31:0] m3s8_addr;
wire  m3s8_cyc;
wire  [31:0] m3s8_data_i;
wire  [31:0] m3s8_data_o;
wire  m3s8_err;
wire  m3s8_rty;
wire  [3:0] m3s8_sel;
wire  m3s8_stb;
wire  m3s8_we;
wire  m3s9_ack;
wire  [31:0] m3s9_addr;
wire  m3s9_cyc;
wire  [31:0] m3s9_data_i;
wire  [31:0] m3s9_data_o;
wire  m3s9_err;
wire  m3s9_rty;
wire  [3:0] m3s9_sel;
wire  m3s9_stb;
wire  m3s9_we;
output  m4_ack_o;
wire  m4_ack_o;
input  [31:0] m4_addr_i;
wire  [31:0] m4_addr_i;
input  m4_cyc_i;
wire  m4_cyc_i;
input  [31:0] m4_data_i;
wire  [31:0] m4_data_i;
output  [31:0] m4_data_o;
wire  [31:0] m4_data_o;
output  m4_err_o;
wire  m4_err_o;
output  m4_rty_o;
wire  m4_rty_o;
input  [3:0] m4_sel_i;
wire  [3:0] m4_sel_i;
input  m4_stb_i;
wire  m4_stb_i;
input  m4_we_i;
wire  m4_we_i;
wire  m4s0_ack;
wire  [31:0] m4s0_addr;
wire  m4s0_cyc;
wire  [31:0] m4s0_data_i;
wire  [31:0] m4s0_data_o;
wire  m4s0_err;
wire  m4s0_rty;
wire  [3:0] m4s0_sel;
wire  m4s0_stb;
wire  m4s0_we;
wire  m4s10_ack;
wire  [31:0] m4s10_addr;
wire  m4s10_cyc;
wire  [31:0] m4s10_data_i;
wire  [31:0] m4s10_data_o;
wire  m4s10_err;
wire  m4s10_rty;
wire  [3:0] m4s10_sel;
wire  m4s10_stb;
wire  m4s10_we;
wire  m4s11_ack;
wire  [31:0] m4s11_addr;
wire  m4s11_cyc;
wire  [31:0] m4s11_data_i;
wire  [31:0] m4s11_data_o;
wire  m4s11_err;
wire  m4s11_rty;
wire  [3:0] m4s11_sel;
wire  m4s11_stb;
wire  m4s11_we;
wire  m4s12_ack;
wire  [31:0] m4s12_addr;
wire  m4s12_cyc;
wire  [31:0] m4s12_data_i;
wire  [31:0] m4s12_data_o;
wire  m4s12_err;
wire  m4s12_rty;
wire  [3:0] m4s12_sel;
wire  m4s12_stb;
wire  m4s12_we;
wire  m4s13_ack;
wire  [31:0] m4s13_addr;
wire  m4s13_cyc;
wire  [31:0] m4s13_data_i;
wire  [31:0] m4s13_data_o;
wire  m4s13_err;
wire  m4s13_rty;
wire  [3:0] m4s13_sel;
wire  m4s13_stb;
wire  m4s13_we;
wire  m4s14_ack;
wire  [31:0] m4s14_addr;
wire  m4s14_cyc;
wire  [31:0] m4s14_data_i;
wire  [31:0] m4s14_data_o;
wire  m4s14_err;
wire  m4s14_rty;
wire  [3:0] m4s14_sel;
wire  m4s14_stb;
wire  m4s14_we;
wire  m4s15_ack;
wire  [31:0] m4s15_addr;
wire  m4s15_cyc;
wire  [31:0] m4s15_data_i;
wire  [31:0] m4s15_data_o;
wire  m4s15_err;
wire  m4s15_rty;
wire  [3:0] m4s15_sel;
wire  m4s15_stb;
wire  m4s15_we;
wire  m4s1_ack;
wire  [31:0] m4s1_addr;
wire  m4s1_cyc;
wire  [31:0] m4s1_data_i;
wire  [31:0] m4s1_data_o;
wire  m4s1_err;
wire  m4s1_rty;
wire  [3:0] m4s1_sel;
wire  m4s1_stb;
wire  m4s1_we;
wire  m4s2_ack;
wire  [31:0] m4s2_addr;
wire  m4s2_cyc;
wire  [31:0] m4s2_data_i;
wire  [31:0] m4s2_data_o;
wire  m4s2_err;
wire  m4s2_rty;
wire  [3:0] m4s2_sel;
wire  m4s2_stb;
wire  m4s2_we;
wire  m4s3_ack;
wire  [31:0] m4s3_addr;
wire  m4s3_cyc;
wire  [31:0] m4s3_data_i;
wire  [31:0] m4s3_data_o;
wire  m4s3_err;
wire  m4s3_rty;
wire  [3:0] m4s3_sel;
wire  m4s3_stb;
wire  m4s3_we;
wire  m4s4_ack;
wire  [31:0] m4s4_addr;
wire  m4s4_cyc;
wire  [31:0] m4s4_data_i;
wire  [31:0] m4s4_data_o;
wire  m4s4_err;
wire  m4s4_rty;
wire  [3:0] m4s4_sel;
wire  m4s4_stb;
wire  m4s4_we;
wire  m4s5_ack;
wire  [31:0] m4s5_addr;
wire  m4s5_cyc;
wire  [31:0] m4s5_data_i;
wire  [31:0] m4s5_data_o;
wire  m4s5_err;
wire  m4s5_rty;
wire  [3:0] m4s5_sel;
wire  m4s5_stb;
wire  m4s5_we;
wire  m4s6_ack;
wire  [31:0] m4s6_addr;
wire  m4s6_cyc;
wire  [31:0] m4s6_data_i;
wire  [31:0] m4s6_data_o;
wire  m4s6_err;
wire  m4s6_rty;
wire  [3:0] m4s6_sel;
wire  m4s6_stb;
wire  m4s6_we;
wire  m4s7_ack;
wire  [31:0] m4s7_addr;
wire  m4s7_cyc;
wire  [31:0] m4s7_data_i;
wire  [31:0] m4s7_data_o;
wire  m4s7_err;
wire  m4s7_rty;
wire  [3:0] m4s7_sel;
wire  m4s7_stb;
wire  m4s7_we;
wire  m4s8_ack;
wire  [31:0] m4s8_addr;
wire  m4s8_cyc;
wire  [31:0] m4s8_data_i;
wire  [31:0] m4s8_data_o;
wire  m4s8_err;
wire  m4s8_rty;
wire  [3:0] m4s8_sel;
wire  m4s8_stb;
wire  m4s8_we;
wire  m4s9_ack;
wire  [31:0] m4s9_addr;
wire  m4s9_cyc;
wire  [31:0] m4s9_data_i;
wire  [31:0] m4s9_data_o;
wire  m4s9_err;
wire  m4s9_rty;
wire  [3:0] m4s9_sel;
wire  m4s9_stb;
wire  m4s9_we;
output  m5_ack_o;
wire  m5_ack_o;
input  [31:0] m5_addr_i;
wire  [31:0] m5_addr_i;
input  m5_cyc_i;
wire  m5_cyc_i;
input  [31:0] m5_data_i;
wire  [31:0] m5_data_i;
output  [31:0] m5_data_o;
wire  [31:0] m5_data_o;
output  m5_err_o;
wire  m5_err_o;
output  m5_rty_o;
wire  m5_rty_o;
input  [3:0] m5_sel_i;
wire  [3:0] m5_sel_i;
input  m5_stb_i;
wire  m5_stb_i;
input  m5_we_i;
wire  m5_we_i;
wire  m5s0_ack;
wire  [31:0] m5s0_addr;
wire  m5s0_cyc;
wire  [31:0] m5s0_data_i;
wire  [31:0] m5s0_data_o;
wire  m5s0_err;
wire  m5s0_rty;
wire  [3:0] m5s0_sel;
wire  m5s0_stb;
wire  m5s0_we;
wire  m5s10_ack;
wire  [31:0] m5s10_addr;
wire  m5s10_cyc;
wire  [31:0] m5s10_data_i;
wire  [31:0] m5s10_data_o;
wire  m5s10_err;
wire  m5s10_rty;
wire  [3:0] m5s10_sel;
wire  m5s10_stb;
wire  m5s10_we;
wire  m5s11_ack;
wire  [31:0] m5s11_addr;
wire  m5s11_cyc;
wire  [31:0] m5s11_data_i;
wire  [31:0] m5s11_data_o;
wire  m5s11_err;
wire  m5s11_rty;
wire  [3:0] m5s11_sel;
wire  m5s11_stb;
wire  m5s11_we;
wire  m5s12_ack;
wire  [31:0] m5s12_addr;
wire  m5s12_cyc;
wire  [31:0] m5s12_data_i;
wire  [31:0] m5s12_data_o;
wire  m5s12_err;
wire  m5s12_rty;
wire  [3:0] m5s12_sel;
wire  m5s12_stb;
wire  m5s12_we;
wire  m5s13_ack;
wire  [31:0] m5s13_addr;
wire  m5s13_cyc;
wire  [31:0] m5s13_data_i;
wire  [31:0] m5s13_data_o;
wire  m5s13_err;
wire  m5s13_rty;
wire  [3:0] m5s13_sel;
wire  m5s13_stb;
wire  m5s13_we;
wire  m5s14_ack;
wire  [31:0] m5s14_addr;
wire  m5s14_cyc;
wire  [31:0] m5s14_data_i;
wire  [31:0] m5s14_data_o;
wire  m5s14_err;
wire  m5s14_rty;
wire  [3:0] m5s14_sel;
wire  m5s14_stb;
wire  m5s14_we;
wire  m5s15_ack;
wire  [31:0] m5s15_addr;
wire  m5s15_cyc;
wire  [31:0] m5s15_data_i;
wire  [31:0] m5s15_data_o;
wire  m5s15_err;
wire  m5s15_rty;
wire  [3:0] m5s15_sel;
wire  m5s15_stb;
wire  m5s15_we;
wire  m5s1_ack;
wire  [31:0] m5s1_addr;
wire  m5s1_cyc;
wire  [31:0] m5s1_data_i;
wire  [31:0] m5s1_data_o;
wire  m5s1_err;
wire  m5s1_rty;
wire  [3:0] m5s1_sel;
wire  m5s1_stb;
wire  m5s1_we;
wire  m5s2_ack;
wire  [31:0] m5s2_addr;
wire  m5s2_cyc;
wire  [31:0] m5s2_data_i;
wire  [31:0] m5s2_data_o;
wire  m5s2_err;
wire  m5s2_rty;
wire  [3:0] m5s2_sel;
wire  m5s2_stb;
wire  m5s2_we;
wire  m5s3_ack;
wire  [31:0] m5s3_addr;
wire  m5s3_cyc;
wire  [31:0] m5s3_data_i;
wire  [31:0] m5s3_data_o;
wire  m5s3_err;
wire  m5s3_rty;
wire  [3:0] m5s3_sel;
wire  m5s3_stb;
wire  m5s3_we;
wire  m5s4_ack;
wire  [31:0] m5s4_addr;
wire  m5s4_cyc;
wire  [31:0] m5s4_data_i;
wire  [31:0] m5s4_data_o;
wire  m5s4_err;
wire  m5s4_rty;
wire  [3:0] m5s4_sel;
wire  m5s4_stb;
wire  m5s4_we;
wire  m5s5_ack;
wire  [31:0] m5s5_addr;
wire  m5s5_cyc;
wire  [31:0] m5s5_data_i;
wire  [31:0] m5s5_data_o;
wire  m5s5_err;
wire  m5s5_rty;
wire  [3:0] m5s5_sel;
wire  m5s5_stb;
wire  m5s5_we;
wire  m5s6_ack;
wire  [31:0] m5s6_addr;
wire  m5s6_cyc;
wire  [31:0] m5s6_data_i;
wire  [31:0] m5s6_data_o;
wire  m5s6_err;
wire  m5s6_rty;
wire  [3:0] m5s6_sel;
wire  m5s6_stb;
wire  m5s6_we;
wire  m5s7_ack;
wire  [31:0] m5s7_addr;
wire  m5s7_cyc;
wire  [31:0] m5s7_data_i;
wire  [31:0] m5s7_data_o;
wire  m5s7_err;
wire  m5s7_rty;
wire  [3:0] m5s7_sel;
wire  m5s7_stb;
wire  m5s7_we;
wire  m5s8_ack;
wire  [31:0] m5s8_addr;
wire  m5s8_cyc;
wire  [31:0] m5s8_data_i;
wire  [31:0] m5s8_data_o;
wire  m5s8_err;
wire  m5s8_rty;
wire  [3:0] m5s8_sel;
wire  m5s8_stb;
wire  m5s8_we;
wire  m5s9_ack;
wire  [31:0] m5s9_addr;
wire  m5s9_cyc;
wire  [31:0] m5s9_data_i;
wire  [31:0] m5s9_data_o;
wire  m5s9_err;
wire  m5s9_rty;
wire  [3:0] m5s9_sel;
wire  m5s9_stb;
wire  m5s9_we;
output  m6_ack_o;
wire  m6_ack_o;
input  [31:0] m6_addr_i;
wire  [31:0] m6_addr_i;
input  m6_cyc_i;
wire  m6_cyc_i;
input  [31:0] m6_data_i;
wire  [31:0] m6_data_i;
output  [31:0] m6_data_o;
wire  [31:0] m6_data_o;
output  m6_err_o;
wire  m6_err_o;
output  m6_rty_o;
wire  m6_rty_o;
input  [3:0] m6_sel_i;
wire  [3:0] m6_sel_i;
input  m6_stb_i;
wire  m6_stb_i;
input  m6_we_i;
wire  m6_we_i;
wire  m6s0_ack;
wire  [31:0] m6s0_addr;
wire  m6s0_cyc;
wire  [31:0] m6s0_data_i;
wire  [31:0] m6s0_data_o;
wire  m6s0_err;
wire  m6s0_rty;
wire  [3:0] m6s0_sel;
wire  m6s0_stb;
wire  m6s0_we;
wire  m6s10_ack;
wire  [31:0] m6s10_addr;
wire  m6s10_cyc;
wire  [31:0] m6s10_data_i;
wire  [31:0] m6s10_data_o;
wire  m6s10_err;
wire  m6s10_rty;
wire  [3:0] m6s10_sel;
wire  m6s10_stb;
wire  m6s10_we;
wire  m6s11_ack;
wire  [31:0] m6s11_addr;
wire  m6s11_cyc;
wire  [31:0] m6s11_data_i;
wire  [31:0] m6s11_data_o;
wire  m6s11_err;
wire  m6s11_rty;
wire  [3:0] m6s11_sel;
wire  m6s11_stb;
wire  m6s11_we;
wire  m6s12_ack;
wire  [31:0] m6s12_addr;
wire  m6s12_cyc;
wire  [31:0] m6s12_data_i;
wire  [31:0] m6s12_data_o;
wire  m6s12_err;
wire  m6s12_rty;
wire  [3:0] m6s12_sel;
wire  m6s12_stb;
wire  m6s12_we;
wire  m6s13_ack;
wire  [31:0] m6s13_addr;
wire  m6s13_cyc;
wire  [31:0] m6s13_data_i;
wire  [31:0] m6s13_data_o;
wire  m6s13_err;
wire  m6s13_rty;
wire  [3:0] m6s13_sel;
wire  m6s13_stb;
wire  m6s13_we;
wire  m6s14_ack;
wire  [31:0] m6s14_addr;
wire  m6s14_cyc;
wire  [31:0] m6s14_data_i;
wire  [31:0] m6s14_data_o;
wire  m6s14_err;
wire  m6s14_rty;
wire  [3:0] m6s14_sel;
wire  m6s14_stb;
wire  m6s14_we;
wire  m6s15_ack;
wire  [31:0] m6s15_addr;
wire  m6s15_cyc;
wire  [31:0] m6s15_data_i;
wire  [31:0] m6s15_data_o;
wire  m6s15_err;
wire  m6s15_rty;
wire  [3:0] m6s15_sel;
wire  m6s15_stb;
wire  m6s15_we;
wire  m6s1_ack;
wire  [31:0] m6s1_addr;
wire  m6s1_cyc;
wire  [31:0] m6s1_data_i;
wire  [31:0] m6s1_data_o;
wire  m6s1_err;
wire  m6s1_rty;
wire  [3:0] m6s1_sel;
wire  m6s1_stb;
wire  m6s1_we;
wire  m6s2_ack;
wire  [31:0] m6s2_addr;
wire  m6s2_cyc;
wire  [31:0] m6s2_data_i;
wire  [31:0] m6s2_data_o;
wire  m6s2_err;
wire  m6s2_rty;
wire  [3:0] m6s2_sel;
wire  m6s2_stb;
wire  m6s2_we;
wire  m6s3_ack;
wire  [31:0] m6s3_addr;
wire  m6s3_cyc;
wire  [31:0] m6s3_data_i;
wire  [31:0] m6s3_data_o;
wire  m6s3_err;
wire  m6s3_rty;
wire  [3:0] m6s3_sel;
wire  m6s3_stb;
wire  m6s3_we;
wire  m6s4_ack;
wire  [31:0] m6s4_addr;
wire  m6s4_cyc;
wire  [31:0] m6s4_data_i;
wire  [31:0] m6s4_data_o;
wire  m6s4_err;
wire  m6s4_rty;
wire  [3:0] m6s4_sel;
wire  m6s4_stb;
wire  m6s4_we;
wire  m6s5_ack;
wire  [31:0] m6s5_addr;
wire  m6s5_cyc;
wire  [31:0] m6s5_data_i;
wire  [31:0] m6s5_data_o;
wire  m6s5_err;
wire  m6s5_rty;
wire  [3:0] m6s5_sel;
wire  m6s5_stb;
wire  m6s5_we;
wire  m6s6_ack;
wire  [31:0] m6s6_addr;
wire  m6s6_cyc;
wire  [31:0] m6s6_data_i;
wire  [31:0] m6s6_data_o;
wire  m6s6_err;
wire  m6s6_rty;
wire  [3:0] m6s6_sel;
wire  m6s6_stb;
wire  m6s6_we;
wire  m6s7_ack;
wire  [31:0] m6s7_addr;
wire  m6s7_cyc;
wire  [31:0] m6s7_data_i;
wire  [31:0] m6s7_data_o;
wire  m6s7_err;
wire  m6s7_rty;
wire  [3:0] m6s7_sel;
wire  m6s7_stb;
wire  m6s7_we;
wire  m6s8_ack;
wire  [31:0] m6s8_addr;
wire  m6s8_cyc;
wire  [31:0] m6s8_data_i;
wire  [31:0] m6s8_data_o;
wire  m6s8_err;
wire  m6s8_rty;
wire  [3:0] m6s8_sel;
wire  m6s8_stb;
wire  m6s8_we;
wire  m6s9_ack;
wire  [31:0] m6s9_addr;
wire  m6s9_cyc;
wire  [31:0] m6s9_data_i;
wire  [31:0] m6s9_data_o;
wire  m6s9_err;
wire  m6s9_rty;
wire  [3:0] m6s9_sel;
wire  m6s9_stb;
wire  m6s9_we;
output  m7_ack_o;
wire  m7_ack_o;
input  [31:0] m7_addr_i;
wire  [31:0] m7_addr_i;
input  m7_cyc_i;
wire  m7_cyc_i;
input  [31:0] m7_data_i;
wire  [31:0] m7_data_i;
output  [31:0] m7_data_o;
wire  [31:0] m7_data_o;
output  m7_err_o;
wire  m7_err_o;
output  m7_rty_o;
wire  m7_rty_o;
input  [3:0] m7_sel_i;
wire  [3:0] m7_sel_i;
input  m7_stb_i;
wire  m7_stb_i;
input  m7_we_i;
wire  m7_we_i;
wire  m7s0_ack;
wire  [31:0] m7s0_addr;
wire  m7s0_cyc;
wire  [31:0] m7s0_data_i;
wire  [31:0] m7s0_data_o;
wire  m7s0_err;
wire  m7s0_rty;
wire  [3:0] m7s0_sel;
wire  m7s0_stb;
wire  m7s0_we;
wire  m7s10_ack;
wire  [31:0] m7s10_addr;
wire  m7s10_cyc;
wire  [31:0] m7s10_data_i;
wire  [31:0] m7s10_data_o;
wire  m7s10_err;
wire  m7s10_rty;
wire  [3:0] m7s10_sel;
wire  m7s10_stb;
wire  m7s10_we;
wire  m7s11_ack;
wire  [31:0] m7s11_addr;
wire  m7s11_cyc;
wire  [31:0] m7s11_data_i;
wire  [31:0] m7s11_data_o;
wire  m7s11_err;
wire  m7s11_rty;
wire  [3:0] m7s11_sel;
wire  m7s11_stb;
wire  m7s11_we;
wire  m7s12_ack;
wire  [31:0] m7s12_addr;
wire  m7s12_cyc;
wire  [31:0] m7s12_data_i;
wire  [31:0] m7s12_data_o;
wire  m7s12_err;
wire  m7s12_rty;
wire  [3:0] m7s12_sel;
wire  m7s12_stb;
wire  m7s12_we;
wire  m7s13_ack;
wire  [31:0] m7s13_addr;
wire  m7s13_cyc;
wire  [31:0] m7s13_data_i;
wire  [31:0] m7s13_data_o;
wire  m7s13_err;
wire  m7s13_rty;
wire  [3:0] m7s13_sel;
wire  m7s13_stb;
wire  m7s13_we;
wire  m7s14_ack;
wire  [31:0] m7s14_addr;
wire  m7s14_cyc;
wire  [31:0] m7s14_data_i;
wire  [31:0] m7s14_data_o;
wire  m7s14_err;
wire  m7s14_rty;
wire  [3:0] m7s14_sel;
wire  m7s14_stb;
wire  m7s14_we;
wire  m7s15_ack;
wire  [31:0] m7s15_addr;
wire  m7s15_cyc;
wire  [31:0] m7s15_data_i;
wire  [31:0] m7s15_data_o;
wire  m7s15_err;
wire  m7s15_rty;
wire  [3:0] m7s15_sel;
wire  m7s15_stb;
wire  m7s15_we;
wire  m7s1_ack;
wire  [31:0] m7s1_addr;
wire  m7s1_cyc;
wire  [31:0] m7s1_data_i;
wire  [31:0] m7s1_data_o;
wire  m7s1_err;
wire  m7s1_rty;
wire  [3:0] m7s1_sel;
wire  m7s1_stb;
wire  m7s1_we;
wire  m7s2_ack;
wire  [31:0] m7s2_addr;
wire  m7s2_cyc;
wire  [31:0] m7s2_data_i;
wire  [31:0] m7s2_data_o;
wire  m7s2_err;
wire  m7s2_rty;
wire  [3:0] m7s2_sel;
wire  m7s2_stb;
wire  m7s2_we;
wire  m7s3_ack;
wire  [31:0] m7s3_addr;
wire  m7s3_cyc;
wire  [31:0] m7s3_data_i;
wire  [31:0] m7s3_data_o;
wire  m7s3_err;
wire  m7s3_rty;
wire  [3:0] m7s3_sel;
wire  m7s3_stb;
wire  m7s3_we;
wire  m7s4_ack;
wire  [31:0] m7s4_addr;
wire  m7s4_cyc;
wire  [31:0] m7s4_data_i;
wire  [31:0] m7s4_data_o;
wire  m7s4_err;
wire  m7s4_rty;
wire  [3:0] m7s4_sel;
wire  m7s4_stb;
wire  m7s4_we;
wire  m7s5_ack;
wire  [31:0] m7s5_addr;
wire  m7s5_cyc;
wire  [31:0] m7s5_data_i;
wire  [31:0] m7s5_data_o;
wire  m7s5_err;
wire  m7s5_rty;
wire  [3:0] m7s5_sel;
wire  m7s5_stb;
wire  m7s5_we;
wire  m7s6_ack;
wire  [31:0] m7s6_addr;
wire  m7s6_cyc;
wire  [31:0] m7s6_data_i;
wire  [31:0] m7s6_data_o;
wire  m7s6_err;
wire  m7s6_rty;
wire  [3:0] m7s6_sel;
wire  m7s6_stb;
wire  m7s6_we;
wire  m7s7_ack;
wire  [31:0] m7s7_addr;
wire  m7s7_cyc;
wire  [31:0] m7s7_data_i;
wire  [31:0] m7s7_data_o;
wire  m7s7_err;
wire  m7s7_rty;
wire  [3:0] m7s7_sel;
wire  m7s7_stb;
wire  m7s7_we;
wire  m7s8_ack;
wire  [31:0] m7s8_addr;
wire  m7s8_cyc;
wire  [31:0] m7s8_data_i;
wire  [31:0] m7s8_data_o;
wire  m7s8_err;
wire  m7s8_rty;
wire  [3:0] m7s8_sel;
wire  m7s8_stb;
wire  m7s8_we;
wire  m7s9_ack;
wire  [31:0] m7s9_addr;
wire  m7s9_cyc;
wire  [31:0] m7s9_data_i;
wire  [31:0] m7s9_data_o;
wire  m7s9_err;
wire  m7s9_rty;
wire  [3:0] m7s9_sel;
wire  m7s9_stb;
wire  m7s9_we;
input  rst_i;
wire  rst_i;
input  s0_ack_i;
wire  s0_ack_i;
output  [31:0] s0_addr_o;
wire  [31:0] s0_addr_o;
output  s0_cyc_o;
wire  s0_cyc_o;
input  [31:0] s0_data_i;
wire  [31:0] s0_data_i;
output  [31:0] s0_data_o;
wire  [31:0] s0_data_o;
input  s0_err_i;
wire  s0_err_i;
input  s0_rty_i;
wire  s0_rty_i;
output  [3:0] s0_sel_o;
wire  [3:0] s0_sel_o;
output  s0_stb_o;
wire  s0_stb_o;
output  s0_we_o;
wire  s0_we_o;
input  s10_ack_i;
wire  s10_ack_i;
output  [31:0] s10_addr_o;
wire  [31:0] s10_addr_o;
output  s10_cyc_o;
wire  s10_cyc_o;
input  [31:0] s10_data_i;
wire  [31:0] s10_data_i;
output  [31:0] s10_data_o;
wire  [31:0] s10_data_o;
input  s10_err_i;
wire  s10_err_i;
input  s10_rty_i;
wire  s10_rty_i;
output  [3:0] s10_sel_o;
wire  [3:0] s10_sel_o;
output  s10_stb_o;
wire  s10_stb_o;
output  s10_we_o;
wire  s10_we_o;
input  s11_ack_i;
wire  s11_ack_i;
output  [31:0] s11_addr_o;
wire  [31:0] s11_addr_o;
output  s11_cyc_o;
wire  s11_cyc_o;
input  [31:0] s11_data_i;
wire  [31:0] s11_data_i;
output  [31:0] s11_data_o;
wire  [31:0] s11_data_o;
input  s11_err_i;
wire  s11_err_i;
input  s11_rty_i;
wire  s11_rty_i;
output  [3:0] s11_sel_o;
wire  [3:0] s11_sel_o;
output  s11_stb_o;
wire  s11_stb_o;
output  s11_we_o;
wire  s11_we_o;
input  s12_ack_i;
wire  s12_ack_i;
output  [31:0] s12_addr_o;
wire  [31:0] s12_addr_o;
output  s12_cyc_o;
wire  s12_cyc_o;
input  [31:0] s12_data_i;
wire  [31:0] s12_data_i;
output  [31:0] s12_data_o;
wire  [31:0] s12_data_o;
input  s12_err_i;
wire  s12_err_i;
input  s12_rty_i;
wire  s12_rty_i;
output  [3:0] s12_sel_o;
wire  [3:0] s12_sel_o;
output  s12_stb_o;
wire  s12_stb_o;
output  s12_we_o;
wire  s12_we_o;
input  s13_ack_i;
wire  s13_ack_i;
output  [31:0] s13_addr_o;
wire  [31:0] s13_addr_o;
output  s13_cyc_o;
wire  s13_cyc_o;
input  [31:0] s13_data_i;
wire  [31:0] s13_data_i;
output  [31:0] s13_data_o;
wire  [31:0] s13_data_o;
input  s13_err_i;
wire  s13_err_i;
input  s13_rty_i;
wire  s13_rty_i;
output  [3:0] s13_sel_o;
wire  [3:0] s13_sel_o;
output  s13_stb_o;
wire  s13_stb_o;
output  s13_we_o;
wire  s13_we_o;
input  s14_ack_i;
wire  s14_ack_i;
output  [31:0] s14_addr_o;
wire  [31:0] s14_addr_o;
output  s14_cyc_o;
wire  s14_cyc_o;
input  [31:0] s14_data_i;
wire  [31:0] s14_data_i;
output  [31:0] s14_data_o;
wire  [31:0] s14_data_o;
input  s14_err_i;
wire  s14_err_i;
input  s14_rty_i;
wire  s14_rty_i;
output  [3:0] s14_sel_o;
wire  [3:0] s14_sel_o;
output  s14_stb_o;
wire  s14_stb_o;
output  s14_we_o;
wire  s14_we_o;
input  s15_ack_i;
wire  s15_ack_i;
output  [31:0] s15_addr_o;
wire  [31:0] s15_addr_o;
output  s15_cyc_o;
wire  s15_cyc_o;
input  [31:0] s15_data_i;
wire  [31:0] s15_data_i;
output  [31:0] s15_data_o;
wire  [31:0] s15_data_o;
input  s15_err_i;
wire  s15_err_i;
input  s15_rty_i;
wire  s15_rty_i;
output  [3:0] s15_sel_o;
wire  [3:0] s15_sel_o;
output  s15_stb_o;
wire  s15_stb_o;
output  s15_we_o;
wire  s15_we_o;
input  s1_ack_i;
wire  s1_ack_i;
output  [31:0] s1_addr_o;
wire  [31:0] s1_addr_o;
output  s1_cyc_o;
wire  s1_cyc_o;
input  [31:0] s1_data_i;
wire  [31:0] s1_data_i;
output  [31:0] s1_data_o;
wire  [31:0] s1_data_o;
input  s1_err_i;
wire  s1_err_i;
input  s1_rty_i;
wire  s1_rty_i;
output  [3:0] s1_sel_o;
wire  [3:0] s1_sel_o;
output  s1_stb_o;
wire  s1_stb_o;
output  s1_we_o;
wire  s1_we_o;
input  s2_ack_i;
wire  s2_ack_i;
output  [31:0] s2_addr_o;
wire  [31:0] s2_addr_o;
output  s2_cyc_o;
wire  s2_cyc_o;
input  [31:0] s2_data_i;
wire  [31:0] s2_data_i;
output  [31:0] s2_data_o;
wire  [31:0] s2_data_o;
input  s2_err_i;
wire  s2_err_i;
input  s2_rty_i;
wire  s2_rty_i;
output  [3:0] s2_sel_o;
wire  [3:0] s2_sel_o;
output  s2_stb_o;
wire  s2_stb_o;
output  s2_we_o;
wire  s2_we_o;
input  s3_ack_i;
wire  s3_ack_i;
output  [31:0] s3_addr_o;
wire  [31:0] s3_addr_o;
output  s3_cyc_o;
wire  s3_cyc_o;
input  [31:0] s3_data_i;
wire  [31:0] s3_data_i;
output  [31:0] s3_data_o;
wire  [31:0] s3_data_o;
input  s3_err_i;
wire  s3_err_i;
input  s3_rty_i;
wire  s3_rty_i;
output  [3:0] s3_sel_o;
wire  [3:0] s3_sel_o;
output  s3_stb_o;
wire  s3_stb_o;
output  s3_we_o;
wire  s3_we_o;
input  s4_ack_i;
wire  s4_ack_i;
output  [31:0] s4_addr_o;
wire  [31:0] s4_addr_o;
output  s4_cyc_o;
wire  s4_cyc_o;
input  [31:0] s4_data_i;
wire  [31:0] s4_data_i;
output  [31:0] s4_data_o;
wire  [31:0] s4_data_o;
input  s4_err_i;
wire  s4_err_i;
input  s4_rty_i;
wire  s4_rty_i;
output  [3:0] s4_sel_o;
wire  [3:0] s4_sel_o;
output  s4_stb_o;
wire  s4_stb_o;
output  s4_we_o;
wire  s4_we_o;
input  s5_ack_i;
wire  s5_ack_i;
output  [31:0] s5_addr_o;
wire  [31:0] s5_addr_o;
output  s5_cyc_o;
wire  s5_cyc_o;
input  [31:0] s5_data_i;
wire  [31:0] s5_data_i;
output  [31:0] s5_data_o;
wire  [31:0] s5_data_o;
input  s5_err_i;
wire  s5_err_i;
input  s5_rty_i;
wire  s5_rty_i;
output  [3:0] s5_sel_o;
wire  [3:0] s5_sel_o;
output  s5_stb_o;
wire  s5_stb_o;
output  s5_we_o;
wire  s5_we_o;
input  s6_ack_i;
wire  s6_ack_i;
output  [31:0] s6_addr_o;
wire  [31:0] s6_addr_o;
output  s6_cyc_o;
wire  s6_cyc_o;
input  [31:0] s6_data_i;
wire  [31:0] s6_data_i;
output  [31:0] s6_data_o;
wire  [31:0] s6_data_o;
input  s6_err_i;
wire  s6_err_i;
input  s6_rty_i;
wire  s6_rty_i;
output  [3:0] s6_sel_o;
wire  [3:0] s6_sel_o;
output  s6_stb_o;
wire  s6_stb_o;
output  s6_we_o;
wire  s6_we_o;
input  s7_ack_i;
wire  s7_ack_i;
output  [31:0] s7_addr_o;
wire  [31:0] s7_addr_o;
output  s7_cyc_o;
wire  s7_cyc_o;
input  [31:0] s7_data_i;
wire  [31:0] s7_data_i;
output  [31:0] s7_data_o;
wire  [31:0] s7_data_o;
input  s7_err_i;
wire  s7_err_i;
input  s7_rty_i;
wire  s7_rty_i;
output  [3:0] s7_sel_o;
wire  [3:0] s7_sel_o;
output  s7_stb_o;
wire  s7_stb_o;
output  s7_we_o;
wire  s7_we_o;
input  s8_ack_i;
wire  s8_ack_i;
output  [31:0] s8_addr_o;
wire  [31:0] s8_addr_o;
output  s8_cyc_o;
wire  s8_cyc_o;
input  [31:0] s8_data_i;
wire  [31:0] s8_data_i;
output  [31:0] s8_data_o;
wire  [31:0] s8_data_o;
input  s8_err_i;
wire  s8_err_i;
input  s8_rty_i;
wire  s8_rty_i;
output  [3:0] s8_sel_o;
wire  [3:0] s8_sel_o;
output  s8_stb_o;
wire  s8_stb_o;
output  s8_we_o;
wire  s8_we_o;
input  s9_ack_i;
wire  s9_ack_i;
output  [31:0] s9_addr_o;
wire  [31:0] s9_addr_o;
output  s9_cyc_o;
wire  s9_cyc_o;
input  [31:0] s9_data_i;
wire  [31:0] s9_data_i;
output  [31:0] s9_data_o;
wire  [31:0] s9_data_o;
input  s9_err_i;
wire  s9_err_i;
input  s9_rty_i;
wire  s9_rty_i;
output  [3:0] s9_sel_o;
wire  [3:0] s9_sel_o;
output  s9_stb_o;
wire  s9_stb_o;
output  s9_we_o;
wire  s9_we_o;
BUFG  _0243_ (
    .I(_0000_),
    .O(_0001_)
  );
IBUF  _0244_ (
    .I(clk_i),
    .O(_0000_)
  );
OBUF  _0245_ (
    .I(_0002_),
    .O(m0_ack_o)
  );
IBUF  _0246_ (
    .I(m0_addr_i[0]),
    .O(_0003_[0])
  );
IBUF  _0247_ (
    .I(m0_addr_i[1]),
    .O(_0003_[1])
  );
IBUF  _0248_ (
    .I(m0_addr_i[10]),
    .O(_0003_[10])
  );
IBUF  _0249_ (
    .I(m0_addr_i[11]),
    .O(_0003_[11])
  );
IBUF  _0250_ (
    .I(m0_addr_i[12]),
    .O(_0003_[12])
  );
IBUF  _0251_ (
    .I(m0_addr_i[13]),
    .O(_0003_[13])
  );
IBUF  _0252_ (
    .I(m0_addr_i[14]),
    .O(_0003_[14])
  );
IBUF  _0253_ (
    .I(m0_addr_i[15]),
    .O(_0003_[15])
  );
IBUF  _0254_ (
    .I(m0_addr_i[16]),
    .O(_0003_[16])
  );
IBUF  _0255_ (
    .I(m0_addr_i[17]),
    .O(_0003_[17])
  );
IBUF  _0256_ (
    .I(m0_addr_i[18]),
    .O(_0003_[18])
  );
IBUF  _0257_ (
    .I(m0_addr_i[19]),
    .O(_0003_[19])
  );
IBUF  _0258_ (
    .I(m0_addr_i[2]),
    .O(_0003_[2])
  );
IBUF  _0259_ (
    .I(m0_addr_i[20]),
    .O(_0003_[20])
  );
IBUF  _0260_ (
    .I(m0_addr_i[21]),
    .O(_0003_[21])
  );
IBUF  _0261_ (
    .I(m0_addr_i[22]),
    .O(_0003_[22])
  );
IBUF  _0262_ (
    .I(m0_addr_i[23]),
    .O(_0003_[23])
  );
IBUF  _0263_ (
    .I(m0_addr_i[24]),
    .O(_0003_[24])
  );
IBUF  _0264_ (
    .I(m0_addr_i[25]),
    .O(_0003_[25])
  );
IBUF  _0265_ (
    .I(m0_addr_i[26]),
    .O(_0003_[26])
  );
IBUF  _0266_ (
    .I(m0_addr_i[27]),
    .O(_0003_[27])
  );
IBUF  _0267_ (
    .I(m0_addr_i[28]),
    .O(_0003_[28])
  );
IBUF  _0268_ (
    .I(m0_addr_i[29]),
    .O(_0003_[29])
  );
IBUF  _0269_ (
    .I(m0_addr_i[3]),
    .O(_0003_[3])
  );
IBUF  _0270_ (
    .I(m0_addr_i[30]),
    .O(_0003_[30])
  );
IBUF  _0271_ (
    .I(m0_addr_i[31]),
    .O(_0003_[31])
  );
IBUF  _0272_ (
    .I(m0_addr_i[4]),
    .O(_0003_[4])
  );
IBUF  _0273_ (
    .I(m0_addr_i[5]),
    .O(_0003_[5])
  );
IBUF  _0274_ (
    .I(m0_addr_i[6]),
    .O(_0003_[6])
  );
IBUF  _0275_ (
    .I(m0_addr_i[7]),
    .O(_0003_[7])
  );
IBUF  _0276_ (
    .I(m0_addr_i[8]),
    .O(_0003_[8])
  );
IBUF  _0277_ (
    .I(m0_addr_i[9]),
    .O(_0003_[9])
  );
IBUF  _0278_ (
    .I(m0_cyc_i),
    .O(_0004_)
  );
IBUF  _0279_ (
    .I(m0_data_i[0]),
    .O(_0005_[0])
  );
IBUF  _0280_ (
    .I(m0_data_i[1]),
    .O(_0005_[1])
  );
IBUF  _0281_ (
    .I(m0_data_i[10]),
    .O(_0005_[10])
  );
IBUF  _0282_ (
    .I(m0_data_i[11]),
    .O(_0005_[11])
  );
IBUF  _0283_ (
    .I(m0_data_i[12]),
    .O(_0005_[12])
  );
IBUF  _0284_ (
    .I(m0_data_i[13]),
    .O(_0005_[13])
  );
IBUF  _0285_ (
    .I(m0_data_i[14]),
    .O(_0005_[14])
  );
IBUF  _0286_ (
    .I(m0_data_i[15]),
    .O(_0005_[15])
  );
IBUF  _0287_ (
    .I(m0_data_i[16]),
    .O(_0005_[16])
  );
IBUF  _0288_ (
    .I(m0_data_i[17]),
    .O(_0005_[17])
  );
IBUF  _0289_ (
    .I(m0_data_i[18]),
    .O(_0005_[18])
  );
IBUF  _0290_ (
    .I(m0_data_i[19]),
    .O(_0005_[19])
  );
IBUF  _0291_ (
    .I(m0_data_i[2]),
    .O(_0005_[2])
  );
IBUF  _0292_ (
    .I(m0_data_i[20]),
    .O(_0005_[20])
  );
IBUF  _0293_ (
    .I(m0_data_i[21]),
    .O(_0005_[21])
  );
IBUF  _0294_ (
    .I(m0_data_i[22]),
    .O(_0005_[22])
  );
IBUF  _0295_ (
    .I(m0_data_i[23]),
    .O(_0005_[23])
  );
IBUF  _0296_ (
    .I(m0_data_i[24]),
    .O(_0005_[24])
  );
IBUF  _0297_ (
    .I(m0_data_i[25]),
    .O(_0005_[25])
  );
IBUF  _0298_ (
    .I(m0_data_i[26]),
    .O(_0005_[26])
  );
IBUF  _0299_ (
    .I(m0_data_i[27]),
    .O(_0005_[27])
  );
IBUF  _0300_ (
    .I(m0_data_i[28]),
    .O(_0005_[28])
  );
IBUF  _0301_ (
    .I(m0_data_i[29]),
    .O(_0005_[29])
  );
IBUF  _0302_ (
    .I(m0_data_i[3]),
    .O(_0005_[3])
  );
IBUF  _0303_ (
    .I(m0_data_i[30]),
    .O(_0005_[30])
  );
IBUF  _0304_ (
    .I(m0_data_i[31]),
    .O(_0005_[31])
  );
IBUF  _0305_ (
    .I(m0_data_i[4]),
    .O(_0005_[4])
  );
IBUF  _0306_ (
    .I(m0_data_i[5]),
    .O(_0005_[5])
  );
IBUF  _0307_ (
    .I(m0_data_i[6]),
    .O(_0005_[6])
  );
IBUF  _0308_ (
    .I(m0_data_i[7]),
    .O(_0005_[7])
  );
IBUF  _0309_ (
    .I(m0_data_i[8]),
    .O(_0005_[8])
  );
IBUF  _0310_ (
    .I(m0_data_i[9]),
    .O(_0005_[9])
  );
OBUF  _0311_ (
    .I(_0006_[0]),
    .O(m0_data_o[0])
  );
OBUF  _0312_ (
    .I(_0006_[1]),
    .O(m0_data_o[1])
  );
OBUF  _0313_ (
    .I(_0006_[10]),
    .O(m0_data_o[10])
  );
OBUF  _0314_ (
    .I(_0006_[11]),
    .O(m0_data_o[11])
  );
OBUF  _0315_ (
    .I(_0006_[12]),
    .O(m0_data_o[12])
  );
OBUF  _0316_ (
    .I(_0006_[13]),
    .O(m0_data_o[13])
  );
OBUF  _0317_ (
    .I(_0006_[14]),
    .O(m0_data_o[14])
  );
OBUF  _0318_ (
    .I(_0006_[15]),
    .O(m0_data_o[15])
  );
OBUF  _0319_ (
    .I(_0006_[16]),
    .O(m0_data_o[16])
  );
OBUF  _0320_ (
    .I(_0006_[17]),
    .O(m0_data_o[17])
  );
OBUF  _0321_ (
    .I(_0006_[18]),
    .O(m0_data_o[18])
  );
OBUF  _0322_ (
    .I(_0006_[19]),
    .O(m0_data_o[19])
  );
OBUF  _0323_ (
    .I(_0006_[2]),
    .O(m0_data_o[2])
  );
OBUF  _0324_ (
    .I(_0006_[20]),
    .O(m0_data_o[20])
  );
OBUF  _0325_ (
    .I(_0006_[21]),
    .O(m0_data_o[21])
  );
OBUF  _0326_ (
    .I(_0006_[22]),
    .O(m0_data_o[22])
  );
OBUF  _0327_ (
    .I(_0006_[23]),
    .O(m0_data_o[23])
  );
OBUF  _0328_ (
    .I(_0006_[24]),
    .O(m0_data_o[24])
  );
OBUF  _0329_ (
    .I(_0006_[25]),
    .O(m0_data_o[25])
  );
OBUF  _0330_ (
    .I(_0006_[26]),
    .O(m0_data_o[26])
  );
OBUF  _0331_ (
    .I(_0006_[27]),
    .O(m0_data_o[27])
  );
OBUF  _0332_ (
    .I(_0006_[28]),
    .O(m0_data_o[28])
  );
OBUF  _0333_ (
    .I(_0006_[29]),
    .O(m0_data_o[29])
  );
OBUF  _0334_ (
    .I(_0006_[3]),
    .O(m0_data_o[3])
  );
OBUF  _0335_ (
    .I(_0006_[30]),
    .O(m0_data_o[30])
  );
OBUF  _0336_ (
    .I(_0006_[31]),
    .O(m0_data_o[31])
  );
OBUF  _0337_ (
    .I(_0006_[4]),
    .O(m0_data_o[4])
  );
OBUF  _0338_ (
    .I(_0006_[5]),
    .O(m0_data_o[5])
  );
OBUF  _0339_ (
    .I(_0006_[6]),
    .O(m0_data_o[6])
  );
OBUF  _0340_ (
    .I(_0006_[7]),
    .O(m0_data_o[7])
  );
OBUF  _0341_ (
    .I(_0006_[8]),
    .O(m0_data_o[8])
  );
OBUF  _0342_ (
    .I(_0006_[9]),
    .O(m0_data_o[9])
  );
OBUF  _0343_ (
    .I(_0007_),
    .O(m0_err_o)
  );
OBUF  _0344_ (
    .I(_0008_),
    .O(m0_rty_o)
  );
IBUF  _0345_ (
    .I(m0_sel_i[0]),
    .O(_0009_[0])
  );
IBUF  _0346_ (
    .I(m0_sel_i[1]),
    .O(_0009_[1])
  );
IBUF  _0347_ (
    .I(m0_sel_i[2]),
    .O(_0009_[2])
  );
IBUF  _0348_ (
    .I(m0_sel_i[3]),
    .O(_0009_[3])
  );
IBUF  _0349_ (
    .I(m0_stb_i),
    .O(_0010_)
  );
IBUF  _0350_ (
    .I(m0_we_i),
    .O(_0011_)
  );
OBUF  _0351_ (
    .I(_0012_),
    .O(m1_ack_o)
  );
IBUF  _0352_ (
    .I(m1_addr_i[0]),
    .O(_0013_[0])
  );
IBUF  _0353_ (
    .I(m1_addr_i[1]),
    .O(_0013_[1])
  );
IBUF  _0354_ (
    .I(m1_addr_i[10]),
    .O(_0013_[10])
  );
IBUF  _0355_ (
    .I(m1_addr_i[11]),
    .O(_0013_[11])
  );
IBUF  _0356_ (
    .I(m1_addr_i[12]),
    .O(_0013_[12])
  );
IBUF  _0357_ (
    .I(m1_addr_i[13]),
    .O(_0013_[13])
  );
IBUF  _0358_ (
    .I(m1_addr_i[14]),
    .O(_0013_[14])
  );
IBUF  _0359_ (
    .I(m1_addr_i[15]),
    .O(_0013_[15])
  );
IBUF  _0360_ (
    .I(m1_addr_i[16]),
    .O(_0013_[16])
  );
IBUF  _0361_ (
    .I(m1_addr_i[17]),
    .O(_0013_[17])
  );
IBUF  _0362_ (
    .I(m1_addr_i[18]),
    .O(_0013_[18])
  );
IBUF  _0363_ (
    .I(m1_addr_i[19]),
    .O(_0013_[19])
  );
IBUF  _0364_ (
    .I(m1_addr_i[2]),
    .O(_0013_[2])
  );
IBUF  _0365_ (
    .I(m1_addr_i[20]),
    .O(_0013_[20])
  );
IBUF  _0366_ (
    .I(m1_addr_i[21]),
    .O(_0013_[21])
  );
IBUF  _0367_ (
    .I(m1_addr_i[22]),
    .O(_0013_[22])
  );
IBUF  _0368_ (
    .I(m1_addr_i[23]),
    .O(_0013_[23])
  );
IBUF  _0369_ (
    .I(m1_addr_i[24]),
    .O(_0013_[24])
  );
IBUF  _0370_ (
    .I(m1_addr_i[25]),
    .O(_0013_[25])
  );
IBUF  _0371_ (
    .I(m1_addr_i[26]),
    .O(_0013_[26])
  );
IBUF  _0372_ (
    .I(m1_addr_i[27]),
    .O(_0013_[27])
  );
IBUF  _0373_ (
    .I(m1_addr_i[28]),
    .O(_0013_[28])
  );
IBUF  _0374_ (
    .I(m1_addr_i[29]),
    .O(_0013_[29])
  );
IBUF  _0375_ (
    .I(m1_addr_i[3]),
    .O(_0013_[3])
  );
IBUF  _0376_ (
    .I(m1_addr_i[30]),
    .O(_0013_[30])
  );
IBUF  _0377_ (
    .I(m1_addr_i[31]),
    .O(_0013_[31])
  );
IBUF  _0378_ (
    .I(m1_addr_i[4]),
    .O(_0013_[4])
  );
IBUF  _0379_ (
    .I(m1_addr_i[5]),
    .O(_0013_[5])
  );
IBUF  _0380_ (
    .I(m1_addr_i[6]),
    .O(_0013_[6])
  );
IBUF  _0381_ (
    .I(m1_addr_i[7]),
    .O(_0013_[7])
  );
IBUF  _0382_ (
    .I(m1_addr_i[8]),
    .O(_0013_[8])
  );
IBUF  _0383_ (
    .I(m1_addr_i[9]),
    .O(_0013_[9])
  );
IBUF  _0384_ (
    .I(m1_cyc_i),
    .O(_0014_)
  );
IBUF  _0385_ (
    .I(m1_data_i[0]),
    .O(_0015_[0])
  );
IBUF  _0386_ (
    .I(m1_data_i[1]),
    .O(_0015_[1])
  );
IBUF  _0387_ (
    .I(m1_data_i[10]),
    .O(_0015_[10])
  );
IBUF  _0388_ (
    .I(m1_data_i[11]),
    .O(_0015_[11])
  );
IBUF  _0389_ (
    .I(m1_data_i[12]),
    .O(_0015_[12])
  );
IBUF  _0390_ (
    .I(m1_data_i[13]),
    .O(_0015_[13])
  );
IBUF  _0391_ (
    .I(m1_data_i[14]),
    .O(_0015_[14])
  );
IBUF  _0392_ (
    .I(m1_data_i[15]),
    .O(_0015_[15])
  );
IBUF  _0393_ (
    .I(m1_data_i[16]),
    .O(_0015_[16])
  );
IBUF  _0394_ (
    .I(m1_data_i[17]),
    .O(_0015_[17])
  );
IBUF  _0395_ (
    .I(m1_data_i[18]),
    .O(_0015_[18])
  );
IBUF  _0396_ (
    .I(m1_data_i[19]),
    .O(_0015_[19])
  );
IBUF  _0397_ (
    .I(m1_data_i[2]),
    .O(_0015_[2])
  );
IBUF  _0398_ (
    .I(m1_data_i[20]),
    .O(_0015_[20])
  );
IBUF  _0399_ (
    .I(m1_data_i[21]),
    .O(_0015_[21])
  );
IBUF  _0400_ (
    .I(m1_data_i[22]),
    .O(_0015_[22])
  );
IBUF  _0401_ (
    .I(m1_data_i[23]),
    .O(_0015_[23])
  );
IBUF  _0402_ (
    .I(m1_data_i[24]),
    .O(_0015_[24])
  );
IBUF  _0403_ (
    .I(m1_data_i[25]),
    .O(_0015_[25])
  );
IBUF  _0404_ (
    .I(m1_data_i[26]),
    .O(_0015_[26])
  );
IBUF  _0405_ (
    .I(m1_data_i[27]),
    .O(_0015_[27])
  );
IBUF  _0406_ (
    .I(m1_data_i[28]),
    .O(_0015_[28])
  );
IBUF  _0407_ (
    .I(m1_data_i[29]),
    .O(_0015_[29])
  );
IBUF  _0408_ (
    .I(m1_data_i[3]),
    .O(_0015_[3])
  );
IBUF  _0409_ (
    .I(m1_data_i[30]),
    .O(_0015_[30])
  );
IBUF  _0410_ (
    .I(m1_data_i[31]),
    .O(_0015_[31])
  );
IBUF  _0411_ (
    .I(m1_data_i[4]),
    .O(_0015_[4])
  );
IBUF  _0412_ (
    .I(m1_data_i[5]),
    .O(_0015_[5])
  );
IBUF  _0413_ (
    .I(m1_data_i[6]),
    .O(_0015_[6])
  );
IBUF  _0414_ (
    .I(m1_data_i[7]),
    .O(_0015_[7])
  );
IBUF  _0415_ (
    .I(m1_data_i[8]),
    .O(_0015_[8])
  );
IBUF  _0416_ (
    .I(m1_data_i[9]),
    .O(_0015_[9])
  );
OBUF  _0417_ (
    .I(_0016_[0]),
    .O(m1_data_o[0])
  );
OBUF  _0418_ (
    .I(_0016_[1]),
    .O(m1_data_o[1])
  );
OBUF  _0419_ (
    .I(_0016_[10]),
    .O(m1_data_o[10])
  );
OBUF  _0420_ (
    .I(_0016_[11]),
    .O(m1_data_o[11])
  );
OBUF  _0421_ (
    .I(_0016_[12]),
    .O(m1_data_o[12])
  );
OBUF  _0422_ (
    .I(_0016_[13]),
    .O(m1_data_o[13])
  );
OBUF  _0423_ (
    .I(_0016_[14]),
    .O(m1_data_o[14])
  );
OBUF  _0424_ (
    .I(_0016_[15]),
    .O(m1_data_o[15])
  );
OBUF  _0425_ (
    .I(_0016_[16]),
    .O(m1_data_o[16])
  );
OBUF  _0426_ (
    .I(_0016_[17]),
    .O(m1_data_o[17])
  );
OBUF  _0427_ (
    .I(_0016_[18]),
    .O(m1_data_o[18])
  );
OBUF  _0428_ (
    .I(_0016_[19]),
    .O(m1_data_o[19])
  );
OBUF  _0429_ (
    .I(_0016_[2]),
    .O(m1_data_o[2])
  );
OBUF  _0430_ (
    .I(_0016_[20]),
    .O(m1_data_o[20])
  );
OBUF  _0431_ (
    .I(_0016_[21]),
    .O(m1_data_o[21])
  );
OBUF  _0432_ (
    .I(_0016_[22]),
    .O(m1_data_o[22])
  );
OBUF  _0433_ (
    .I(_0016_[23]),
    .O(m1_data_o[23])
  );
OBUF  _0434_ (
    .I(_0016_[24]),
    .O(m1_data_o[24])
  );
OBUF  _0435_ (
    .I(_0016_[25]),
    .O(m1_data_o[25])
  );
OBUF  _0436_ (
    .I(_0016_[26]),
    .O(m1_data_o[26])
  );
OBUF  _0437_ (
    .I(_0016_[27]),
    .O(m1_data_o[27])
  );
OBUF  _0438_ (
    .I(_0016_[28]),
    .O(m1_data_o[28])
  );
OBUF  _0439_ (
    .I(_0016_[29]),
    .O(m1_data_o[29])
  );
OBUF  _0440_ (
    .I(_0016_[3]),
    .O(m1_data_o[3])
  );
OBUF  _0441_ (
    .I(_0016_[30]),
    .O(m1_data_o[30])
  );
OBUF  _0442_ (
    .I(_0016_[31]),
    .O(m1_data_o[31])
  );
OBUF  _0443_ (
    .I(_0016_[4]),
    .O(m1_data_o[4])
  );
OBUF  _0444_ (
    .I(_0016_[5]),
    .O(m1_data_o[5])
  );
OBUF  _0445_ (
    .I(_0016_[6]),
    .O(m1_data_o[6])
  );
OBUF  _0446_ (
    .I(_0016_[7]),
    .O(m1_data_o[7])
  );
OBUF  _0447_ (
    .I(_0016_[8]),
    .O(m1_data_o[8])
  );
OBUF  _0448_ (
    .I(_0016_[9]),
    .O(m1_data_o[9])
  );
OBUF  _0449_ (
    .I(_0017_),
    .O(m1_err_o)
  );
OBUF  _0450_ (
    .I(_0018_),
    .O(m1_rty_o)
  );
IBUF  _0451_ (
    .I(m1_sel_i[0]),
    .O(_0019_[0])
  );
IBUF  _0452_ (
    .I(m1_sel_i[1]),
    .O(_0019_[1])
  );
IBUF  _0453_ (
    .I(m1_sel_i[2]),
    .O(_0019_[2])
  );
IBUF  _0454_ (
    .I(m1_sel_i[3]),
    .O(_0019_[3])
  );
IBUF  _0455_ (
    .I(m1_stb_i),
    .O(_0020_)
  );
IBUF  _0456_ (
    .I(m1_we_i),
    .O(_0021_)
  );
OBUF  _0457_ (
    .I(_0022_),
    .O(m2_ack_o)
  );
IBUF  _0458_ (
    .I(m2_addr_i[0]),
    .O(_0023_[0])
  );
IBUF  _0459_ (
    .I(m2_addr_i[1]),
    .O(_0023_[1])
  );
IBUF  _0460_ (
    .I(m2_addr_i[10]),
    .O(_0023_[10])
  );
IBUF  _0461_ (
    .I(m2_addr_i[11]),
    .O(_0023_[11])
  );
IBUF  _0462_ (
    .I(m2_addr_i[12]),
    .O(_0023_[12])
  );
IBUF  _0463_ (
    .I(m2_addr_i[13]),
    .O(_0023_[13])
  );
IBUF  _0464_ (
    .I(m2_addr_i[14]),
    .O(_0023_[14])
  );
IBUF  _0465_ (
    .I(m2_addr_i[15]),
    .O(_0023_[15])
  );
IBUF  _0466_ (
    .I(m2_addr_i[16]),
    .O(_0023_[16])
  );
IBUF  _0467_ (
    .I(m2_addr_i[17]),
    .O(_0023_[17])
  );
IBUF  _0468_ (
    .I(m2_addr_i[18]),
    .O(_0023_[18])
  );
IBUF  _0469_ (
    .I(m2_addr_i[19]),
    .O(_0023_[19])
  );
IBUF  _0470_ (
    .I(m2_addr_i[2]),
    .O(_0023_[2])
  );
IBUF  _0471_ (
    .I(m2_addr_i[20]),
    .O(_0023_[20])
  );
IBUF  _0472_ (
    .I(m2_addr_i[21]),
    .O(_0023_[21])
  );
IBUF  _0473_ (
    .I(m2_addr_i[22]),
    .O(_0023_[22])
  );
IBUF  _0474_ (
    .I(m2_addr_i[23]),
    .O(_0023_[23])
  );
IBUF  _0475_ (
    .I(m2_addr_i[24]),
    .O(_0023_[24])
  );
IBUF  _0476_ (
    .I(m2_addr_i[25]),
    .O(_0023_[25])
  );
IBUF  _0477_ (
    .I(m2_addr_i[26]),
    .O(_0023_[26])
  );
IBUF  _0478_ (
    .I(m2_addr_i[27]),
    .O(_0023_[27])
  );
IBUF  _0479_ (
    .I(m2_addr_i[28]),
    .O(_0023_[28])
  );
IBUF  _0480_ (
    .I(m2_addr_i[29]),
    .O(_0023_[29])
  );
IBUF  _0481_ (
    .I(m2_addr_i[3]),
    .O(_0023_[3])
  );
IBUF  _0482_ (
    .I(m2_addr_i[30]),
    .O(_0023_[30])
  );
IBUF  _0483_ (
    .I(m2_addr_i[31]),
    .O(_0023_[31])
  );
IBUF  _0484_ (
    .I(m2_addr_i[4]),
    .O(_0023_[4])
  );
IBUF  _0485_ (
    .I(m2_addr_i[5]),
    .O(_0023_[5])
  );
IBUF  _0486_ (
    .I(m2_addr_i[6]),
    .O(_0023_[6])
  );
IBUF  _0487_ (
    .I(m2_addr_i[7]),
    .O(_0023_[7])
  );
IBUF  _0488_ (
    .I(m2_addr_i[8]),
    .O(_0023_[8])
  );
IBUF  _0489_ (
    .I(m2_addr_i[9]),
    .O(_0023_[9])
  );
IBUF  _0490_ (
    .I(m2_cyc_i),
    .O(_0024_)
  );
IBUF  _0491_ (
    .I(m2_data_i[0]),
    .O(_0025_[0])
  );
IBUF  _0492_ (
    .I(m2_data_i[1]),
    .O(_0025_[1])
  );
IBUF  _0493_ (
    .I(m2_data_i[10]),
    .O(_0025_[10])
  );
IBUF  _0494_ (
    .I(m2_data_i[11]),
    .O(_0025_[11])
  );
IBUF  _0495_ (
    .I(m2_data_i[12]),
    .O(_0025_[12])
  );
IBUF  _0496_ (
    .I(m2_data_i[13]),
    .O(_0025_[13])
  );
IBUF  _0497_ (
    .I(m2_data_i[14]),
    .O(_0025_[14])
  );
IBUF  _0498_ (
    .I(m2_data_i[15]),
    .O(_0025_[15])
  );
IBUF  _0499_ (
    .I(m2_data_i[16]),
    .O(_0025_[16])
  );
IBUF  _0500_ (
    .I(m2_data_i[17]),
    .O(_0025_[17])
  );
IBUF  _0501_ (
    .I(m2_data_i[18]),
    .O(_0025_[18])
  );
IBUF  _0502_ (
    .I(m2_data_i[19]),
    .O(_0025_[19])
  );
IBUF  _0503_ (
    .I(m2_data_i[2]),
    .O(_0025_[2])
  );
IBUF  _0504_ (
    .I(m2_data_i[20]),
    .O(_0025_[20])
  );
IBUF  _0505_ (
    .I(m2_data_i[21]),
    .O(_0025_[21])
  );
IBUF  _0506_ (
    .I(m2_data_i[22]),
    .O(_0025_[22])
  );
IBUF  _0507_ (
    .I(m2_data_i[23]),
    .O(_0025_[23])
  );
IBUF  _0508_ (
    .I(m2_data_i[24]),
    .O(_0025_[24])
  );
IBUF  _0509_ (
    .I(m2_data_i[25]),
    .O(_0025_[25])
  );
IBUF  _0510_ (
    .I(m2_data_i[26]),
    .O(_0025_[26])
  );
IBUF  _0511_ (
    .I(m2_data_i[27]),
    .O(_0025_[27])
  );
IBUF  _0512_ (
    .I(m2_data_i[28]),
    .O(_0025_[28])
  );
IBUF  _0513_ (
    .I(m2_data_i[29]),
    .O(_0025_[29])
  );
IBUF  _0514_ (
    .I(m2_data_i[3]),
    .O(_0025_[3])
  );
IBUF  _0515_ (
    .I(m2_data_i[30]),
    .O(_0025_[30])
  );
IBUF  _0516_ (
    .I(m2_data_i[31]),
    .O(_0025_[31])
  );
IBUF  _0517_ (
    .I(m2_data_i[4]),
    .O(_0025_[4])
  );
IBUF  _0518_ (
    .I(m2_data_i[5]),
    .O(_0025_[5])
  );
IBUF  _0519_ (
    .I(m2_data_i[6]),
    .O(_0025_[6])
  );
IBUF  _0520_ (
    .I(m2_data_i[7]),
    .O(_0025_[7])
  );
IBUF  _0521_ (
    .I(m2_data_i[8]),
    .O(_0025_[8])
  );
IBUF  _0522_ (
    .I(m2_data_i[9]),
    .O(_0025_[9])
  );
OBUF  _0523_ (
    .I(_0026_[0]),
    .O(m2_data_o[0])
  );
OBUF  _0524_ (
    .I(_0026_[1]),
    .O(m2_data_o[1])
  );
OBUF  _0525_ (
    .I(_0026_[10]),
    .O(m2_data_o[10])
  );
OBUF  _0526_ (
    .I(_0026_[11]),
    .O(m2_data_o[11])
  );
OBUF  _0527_ (
    .I(_0026_[12]),
    .O(m2_data_o[12])
  );
OBUF  _0528_ (
    .I(_0026_[13]),
    .O(m2_data_o[13])
  );
OBUF  _0529_ (
    .I(_0026_[14]),
    .O(m2_data_o[14])
  );
OBUF  _0530_ (
    .I(_0026_[15]),
    .O(m2_data_o[15])
  );
OBUF  _0531_ (
    .I(_0026_[16]),
    .O(m2_data_o[16])
  );
OBUF  _0532_ (
    .I(_0026_[17]),
    .O(m2_data_o[17])
  );
OBUF  _0533_ (
    .I(_0026_[18]),
    .O(m2_data_o[18])
  );
OBUF  _0534_ (
    .I(_0026_[19]),
    .O(m2_data_o[19])
  );
OBUF  _0535_ (
    .I(_0026_[2]),
    .O(m2_data_o[2])
  );
OBUF  _0536_ (
    .I(_0026_[20]),
    .O(m2_data_o[20])
  );
OBUF  _0537_ (
    .I(_0026_[21]),
    .O(m2_data_o[21])
  );
OBUF  _0538_ (
    .I(_0026_[22]),
    .O(m2_data_o[22])
  );
OBUF  _0539_ (
    .I(_0026_[23]),
    .O(m2_data_o[23])
  );
OBUF  _0540_ (
    .I(_0026_[24]),
    .O(m2_data_o[24])
  );
OBUF  _0541_ (
    .I(_0026_[25]),
    .O(m2_data_o[25])
  );
OBUF  _0542_ (
    .I(_0026_[26]),
    .O(m2_data_o[26])
  );
OBUF  _0543_ (
    .I(_0026_[27]),
    .O(m2_data_o[27])
  );
OBUF  _0544_ (
    .I(_0026_[28]),
    .O(m2_data_o[28])
  );
OBUF  _0545_ (
    .I(_0026_[29]),
    .O(m2_data_o[29])
  );
OBUF  _0546_ (
    .I(_0026_[3]),
    .O(m2_data_o[3])
  );
OBUF  _0547_ (
    .I(_0026_[30]),
    .O(m2_data_o[30])
  );
OBUF  _0548_ (
    .I(_0026_[31]),
    .O(m2_data_o[31])
  );
OBUF  _0549_ (
    .I(_0026_[4]),
    .O(m2_data_o[4])
  );
OBUF  _0550_ (
    .I(_0026_[5]),
    .O(m2_data_o[5])
  );
OBUF  _0551_ (
    .I(_0026_[6]),
    .O(m2_data_o[6])
  );
OBUF  _0552_ (
    .I(_0026_[7]),
    .O(m2_data_o[7])
  );
OBUF  _0553_ (
    .I(_0026_[8]),
    .O(m2_data_o[8])
  );
OBUF  _0554_ (
    .I(_0026_[9]),
    .O(m2_data_o[9])
  );
OBUF  _0555_ (
    .I(_0027_),
    .O(m2_err_o)
  );
OBUF  _0556_ (
    .I(_0028_),
    .O(m2_rty_o)
  );
IBUF  _0557_ (
    .I(m2_sel_i[0]),
    .O(_0029_[0])
  );
IBUF  _0558_ (
    .I(m2_sel_i[1]),
    .O(_0029_[1])
  );
IBUF  _0559_ (
    .I(m2_sel_i[2]),
    .O(_0029_[2])
  );
IBUF  _0560_ (
    .I(m2_sel_i[3]),
    .O(_0029_[3])
  );
IBUF  _0561_ (
    .I(m2_stb_i),
    .O(_0030_)
  );
IBUF  _0562_ (
    .I(m2_we_i),
    .O(_0031_)
  );
OBUF  _0563_ (
    .I(_0032_),
    .O(m3_ack_o)
  );
IBUF  _0564_ (
    .I(m3_addr_i[0]),
    .O(_0033_[0])
  );
IBUF  _0565_ (
    .I(m3_addr_i[1]),
    .O(_0033_[1])
  );
IBUF  _0566_ (
    .I(m3_addr_i[10]),
    .O(_0033_[10])
  );
IBUF  _0567_ (
    .I(m3_addr_i[11]),
    .O(_0033_[11])
  );
IBUF  _0568_ (
    .I(m3_addr_i[12]),
    .O(_0033_[12])
  );
IBUF  _0569_ (
    .I(m3_addr_i[13]),
    .O(_0033_[13])
  );
IBUF  _0570_ (
    .I(m3_addr_i[14]),
    .O(_0033_[14])
  );
IBUF  _0571_ (
    .I(m3_addr_i[15]),
    .O(_0033_[15])
  );
IBUF  _0572_ (
    .I(m3_addr_i[16]),
    .O(_0033_[16])
  );
IBUF  _0573_ (
    .I(m3_addr_i[17]),
    .O(_0033_[17])
  );
IBUF  _0574_ (
    .I(m3_addr_i[18]),
    .O(_0033_[18])
  );
IBUF  _0575_ (
    .I(m3_addr_i[19]),
    .O(_0033_[19])
  );
IBUF  _0576_ (
    .I(m3_addr_i[2]),
    .O(_0033_[2])
  );
IBUF  _0577_ (
    .I(m3_addr_i[20]),
    .O(_0033_[20])
  );
IBUF  _0578_ (
    .I(m3_addr_i[21]),
    .O(_0033_[21])
  );
IBUF  _0579_ (
    .I(m3_addr_i[22]),
    .O(_0033_[22])
  );
IBUF  _0580_ (
    .I(m3_addr_i[23]),
    .O(_0033_[23])
  );
IBUF  _0581_ (
    .I(m3_addr_i[24]),
    .O(_0033_[24])
  );
IBUF  _0582_ (
    .I(m3_addr_i[25]),
    .O(_0033_[25])
  );
IBUF  _0583_ (
    .I(m3_addr_i[26]),
    .O(_0033_[26])
  );
IBUF  _0584_ (
    .I(m3_addr_i[27]),
    .O(_0033_[27])
  );
IBUF  _0585_ (
    .I(m3_addr_i[28]),
    .O(_0033_[28])
  );
IBUF  _0586_ (
    .I(m3_addr_i[29]),
    .O(_0033_[29])
  );
IBUF  _0587_ (
    .I(m3_addr_i[3]),
    .O(_0033_[3])
  );
IBUF  _0588_ (
    .I(m3_addr_i[30]),
    .O(_0033_[30])
  );
IBUF  _0589_ (
    .I(m3_addr_i[31]),
    .O(_0033_[31])
  );
IBUF  _0590_ (
    .I(m3_addr_i[4]),
    .O(_0033_[4])
  );
IBUF  _0591_ (
    .I(m3_addr_i[5]),
    .O(_0033_[5])
  );
IBUF  _0592_ (
    .I(m3_addr_i[6]),
    .O(_0033_[6])
  );
IBUF  _0593_ (
    .I(m3_addr_i[7]),
    .O(_0033_[7])
  );
IBUF  _0594_ (
    .I(m3_addr_i[8]),
    .O(_0033_[8])
  );
IBUF  _0595_ (
    .I(m3_addr_i[9]),
    .O(_0033_[9])
  );
IBUF  _0596_ (
    .I(m3_cyc_i),
    .O(_0034_)
  );
IBUF  _0597_ (
    .I(m3_data_i[0]),
    .O(_0035_[0])
  );
IBUF  _0598_ (
    .I(m3_data_i[1]),
    .O(_0035_[1])
  );
IBUF  _0599_ (
    .I(m3_data_i[10]),
    .O(_0035_[10])
  );
IBUF  _0600_ (
    .I(m3_data_i[11]),
    .O(_0035_[11])
  );
IBUF  _0601_ (
    .I(m3_data_i[12]),
    .O(_0035_[12])
  );
IBUF  _0602_ (
    .I(m3_data_i[13]),
    .O(_0035_[13])
  );
IBUF  _0603_ (
    .I(m3_data_i[14]),
    .O(_0035_[14])
  );
IBUF  _0604_ (
    .I(m3_data_i[15]),
    .O(_0035_[15])
  );
IBUF  _0605_ (
    .I(m3_data_i[16]),
    .O(_0035_[16])
  );
IBUF  _0606_ (
    .I(m3_data_i[17]),
    .O(_0035_[17])
  );
IBUF  _0607_ (
    .I(m3_data_i[18]),
    .O(_0035_[18])
  );
IBUF  _0608_ (
    .I(m3_data_i[19]),
    .O(_0035_[19])
  );
IBUF  _0609_ (
    .I(m3_data_i[2]),
    .O(_0035_[2])
  );
IBUF  _0610_ (
    .I(m3_data_i[20]),
    .O(_0035_[20])
  );
IBUF  _0611_ (
    .I(m3_data_i[21]),
    .O(_0035_[21])
  );
IBUF  _0612_ (
    .I(m3_data_i[22]),
    .O(_0035_[22])
  );
IBUF  _0613_ (
    .I(m3_data_i[23]),
    .O(_0035_[23])
  );
IBUF  _0614_ (
    .I(m3_data_i[24]),
    .O(_0035_[24])
  );
IBUF  _0615_ (
    .I(m3_data_i[25]),
    .O(_0035_[25])
  );
IBUF  _0616_ (
    .I(m3_data_i[26]),
    .O(_0035_[26])
  );
IBUF  _0617_ (
    .I(m3_data_i[27]),
    .O(_0035_[27])
  );
IBUF  _0618_ (
    .I(m3_data_i[28]),
    .O(_0035_[28])
  );
IBUF  _0619_ (
    .I(m3_data_i[29]),
    .O(_0035_[29])
  );
IBUF  _0620_ (
    .I(m3_data_i[3]),
    .O(_0035_[3])
  );
IBUF  _0621_ (
    .I(m3_data_i[30]),
    .O(_0035_[30])
  );
IBUF  _0622_ (
    .I(m3_data_i[31]),
    .O(_0035_[31])
  );
IBUF  _0623_ (
    .I(m3_data_i[4]),
    .O(_0035_[4])
  );
IBUF  _0624_ (
    .I(m3_data_i[5]),
    .O(_0035_[5])
  );
IBUF  _0625_ (
    .I(m3_data_i[6]),
    .O(_0035_[6])
  );
IBUF  _0626_ (
    .I(m3_data_i[7]),
    .O(_0035_[7])
  );
IBUF  _0627_ (
    .I(m3_data_i[8]),
    .O(_0035_[8])
  );
IBUF  _0628_ (
    .I(m3_data_i[9]),
    .O(_0035_[9])
  );
OBUF  _0629_ (
    .I(_0036_[0]),
    .O(m3_data_o[0])
  );
OBUF  _0630_ (
    .I(_0036_[1]),
    .O(m3_data_o[1])
  );
OBUF  _0631_ (
    .I(_0036_[10]),
    .O(m3_data_o[10])
  );
OBUF  _0632_ (
    .I(_0036_[11]),
    .O(m3_data_o[11])
  );
OBUF  _0633_ (
    .I(_0036_[12]),
    .O(m3_data_o[12])
  );
OBUF  _0634_ (
    .I(_0036_[13]),
    .O(m3_data_o[13])
  );
OBUF  _0635_ (
    .I(_0036_[14]),
    .O(m3_data_o[14])
  );
OBUF  _0636_ (
    .I(_0036_[15]),
    .O(m3_data_o[15])
  );
OBUF  _0637_ (
    .I(_0036_[16]),
    .O(m3_data_o[16])
  );
OBUF  _0638_ (
    .I(_0036_[17]),
    .O(m3_data_o[17])
  );
OBUF  _0639_ (
    .I(_0036_[18]),
    .O(m3_data_o[18])
  );
OBUF  _0640_ (
    .I(_0036_[19]),
    .O(m3_data_o[19])
  );
OBUF  _0641_ (
    .I(_0036_[2]),
    .O(m3_data_o[2])
  );
OBUF  _0642_ (
    .I(_0036_[20]),
    .O(m3_data_o[20])
  );
OBUF  _0643_ (
    .I(_0036_[21]),
    .O(m3_data_o[21])
  );
OBUF  _0644_ (
    .I(_0036_[22]),
    .O(m3_data_o[22])
  );
OBUF  _0645_ (
    .I(_0036_[23]),
    .O(m3_data_o[23])
  );
OBUF  _0646_ (
    .I(_0036_[24]),
    .O(m3_data_o[24])
  );
OBUF  _0647_ (
    .I(_0036_[25]),
    .O(m3_data_o[25])
  );
OBUF  _0648_ (
    .I(_0036_[26]),
    .O(m3_data_o[26])
  );
OBUF  _0649_ (
    .I(_0036_[27]),
    .O(m3_data_o[27])
  );
OBUF  _0650_ (
    .I(_0036_[28]),
    .O(m3_data_o[28])
  );
OBUF  _0651_ (
    .I(_0036_[29]),
    .O(m3_data_o[29])
  );
OBUF  _0652_ (
    .I(_0036_[3]),
    .O(m3_data_o[3])
  );
OBUF  _0653_ (
    .I(_0036_[30]),
    .O(m3_data_o[30])
  );
OBUF  _0654_ (
    .I(_0036_[31]),
    .O(m3_data_o[31])
  );
OBUF  _0655_ (
    .I(_0036_[4]),
    .O(m3_data_o[4])
  );
OBUF  _0656_ (
    .I(_0036_[5]),
    .O(m3_data_o[5])
  );
OBUF  _0657_ (
    .I(_0036_[6]),
    .O(m3_data_o[6])
  );
OBUF  _0658_ (
    .I(_0036_[7]),
    .O(m3_data_o[7])
  );
OBUF  _0659_ (
    .I(_0036_[8]),
    .O(m3_data_o[8])
  );
OBUF  _0660_ (
    .I(_0036_[9]),
    .O(m3_data_o[9])
  );
OBUF  _0661_ (
    .I(_0037_),
    .O(m3_err_o)
  );
OBUF  _0662_ (
    .I(_0038_),
    .O(m3_rty_o)
  );
IBUF  _0663_ (
    .I(m3_sel_i[0]),
    .O(_0039_[0])
  );
IBUF  _0664_ (
    .I(m3_sel_i[1]),
    .O(_0039_[1])
  );
IBUF  _0665_ (
    .I(m3_sel_i[2]),
    .O(_0039_[2])
  );
IBUF  _0666_ (
    .I(m3_sel_i[3]),
    .O(_0039_[3])
  );
IBUF  _0667_ (
    .I(m3_stb_i),
    .O(_0040_)
  );
IBUF  _0668_ (
    .I(m3_we_i),
    .O(_0041_)
  );
OBUF  _0669_ (
    .I(_0042_),
    .O(m4_ack_o)
  );
IBUF  _0670_ (
    .I(m4_addr_i[0]),
    .O(_0043_[0])
  );
IBUF  _0671_ (
    .I(m4_addr_i[1]),
    .O(_0043_[1])
  );
IBUF  _0672_ (
    .I(m4_addr_i[10]),
    .O(_0043_[10])
  );
IBUF  _0673_ (
    .I(m4_addr_i[11]),
    .O(_0043_[11])
  );
IBUF  _0674_ (
    .I(m4_addr_i[12]),
    .O(_0043_[12])
  );
IBUF  _0675_ (
    .I(m4_addr_i[13]),
    .O(_0043_[13])
  );
IBUF  _0676_ (
    .I(m4_addr_i[14]),
    .O(_0043_[14])
  );
IBUF  _0677_ (
    .I(m4_addr_i[15]),
    .O(_0043_[15])
  );
IBUF  _0678_ (
    .I(m4_addr_i[16]),
    .O(_0043_[16])
  );
IBUF  _0679_ (
    .I(m4_addr_i[17]),
    .O(_0043_[17])
  );
IBUF  _0680_ (
    .I(m4_addr_i[18]),
    .O(_0043_[18])
  );
IBUF  _0681_ (
    .I(m4_addr_i[19]),
    .O(_0043_[19])
  );
IBUF  _0682_ (
    .I(m4_addr_i[2]),
    .O(_0043_[2])
  );
IBUF  _0683_ (
    .I(m4_addr_i[20]),
    .O(_0043_[20])
  );
IBUF  _0684_ (
    .I(m4_addr_i[21]),
    .O(_0043_[21])
  );
IBUF  _0685_ (
    .I(m4_addr_i[22]),
    .O(_0043_[22])
  );
IBUF  _0686_ (
    .I(m4_addr_i[23]),
    .O(_0043_[23])
  );
IBUF  _0687_ (
    .I(m4_addr_i[24]),
    .O(_0043_[24])
  );
IBUF  _0688_ (
    .I(m4_addr_i[25]),
    .O(_0043_[25])
  );
IBUF  _0689_ (
    .I(m4_addr_i[26]),
    .O(_0043_[26])
  );
IBUF  _0690_ (
    .I(m4_addr_i[27]),
    .O(_0043_[27])
  );
IBUF  _0691_ (
    .I(m4_addr_i[28]),
    .O(_0043_[28])
  );
IBUF  _0692_ (
    .I(m4_addr_i[29]),
    .O(_0043_[29])
  );
IBUF  _0693_ (
    .I(m4_addr_i[3]),
    .O(_0043_[3])
  );
IBUF  _0694_ (
    .I(m4_addr_i[30]),
    .O(_0043_[30])
  );
IBUF  _0695_ (
    .I(m4_addr_i[31]),
    .O(_0043_[31])
  );
IBUF  _0696_ (
    .I(m4_addr_i[4]),
    .O(_0043_[4])
  );
IBUF  _0697_ (
    .I(m4_addr_i[5]),
    .O(_0043_[5])
  );
IBUF  _0698_ (
    .I(m4_addr_i[6]),
    .O(_0043_[6])
  );
IBUF  _0699_ (
    .I(m4_addr_i[7]),
    .O(_0043_[7])
  );
IBUF  _0700_ (
    .I(m4_addr_i[8]),
    .O(_0043_[8])
  );
IBUF  _0701_ (
    .I(m4_addr_i[9]),
    .O(_0043_[9])
  );
IBUF  _0702_ (
    .I(m4_cyc_i),
    .O(_0044_)
  );
IBUF  _0703_ (
    .I(m4_data_i[0]),
    .O(_0045_[0])
  );
IBUF  _0704_ (
    .I(m4_data_i[1]),
    .O(_0045_[1])
  );
IBUF  _0705_ (
    .I(m4_data_i[10]),
    .O(_0045_[10])
  );
IBUF  _0706_ (
    .I(m4_data_i[11]),
    .O(_0045_[11])
  );
IBUF  _0707_ (
    .I(m4_data_i[12]),
    .O(_0045_[12])
  );
IBUF  _0708_ (
    .I(m4_data_i[13]),
    .O(_0045_[13])
  );
IBUF  _0709_ (
    .I(m4_data_i[14]),
    .O(_0045_[14])
  );
IBUF  _0710_ (
    .I(m4_data_i[15]),
    .O(_0045_[15])
  );
IBUF  _0711_ (
    .I(m4_data_i[16]),
    .O(_0045_[16])
  );
IBUF  _0712_ (
    .I(m4_data_i[17]),
    .O(_0045_[17])
  );
IBUF  _0713_ (
    .I(m4_data_i[18]),
    .O(_0045_[18])
  );
IBUF  _0714_ (
    .I(m4_data_i[19]),
    .O(_0045_[19])
  );
IBUF  _0715_ (
    .I(m4_data_i[2]),
    .O(_0045_[2])
  );
IBUF  _0716_ (
    .I(m4_data_i[20]),
    .O(_0045_[20])
  );
IBUF  _0717_ (
    .I(m4_data_i[21]),
    .O(_0045_[21])
  );
IBUF  _0718_ (
    .I(m4_data_i[22]),
    .O(_0045_[22])
  );
IBUF  _0719_ (
    .I(m4_data_i[23]),
    .O(_0045_[23])
  );
IBUF  _0720_ (
    .I(m4_data_i[24]),
    .O(_0045_[24])
  );
IBUF  _0721_ (
    .I(m4_data_i[25]),
    .O(_0045_[25])
  );
IBUF  _0722_ (
    .I(m4_data_i[26]),
    .O(_0045_[26])
  );
IBUF  _0723_ (
    .I(m4_data_i[27]),
    .O(_0045_[27])
  );
IBUF  _0724_ (
    .I(m4_data_i[28]),
    .O(_0045_[28])
  );
IBUF  _0725_ (
    .I(m4_data_i[29]),
    .O(_0045_[29])
  );
IBUF  _0726_ (
    .I(m4_data_i[3]),
    .O(_0045_[3])
  );
IBUF  _0727_ (
    .I(m4_data_i[30]),
    .O(_0045_[30])
  );
IBUF  _0728_ (
    .I(m4_data_i[31]),
    .O(_0045_[31])
  );
IBUF  _0729_ (
    .I(m4_data_i[4]),
    .O(_0045_[4])
  );
IBUF  _0730_ (
    .I(m4_data_i[5]),
    .O(_0045_[5])
  );
IBUF  _0731_ (
    .I(m4_data_i[6]),
    .O(_0045_[6])
  );
IBUF  _0732_ (
    .I(m4_data_i[7]),
    .O(_0045_[7])
  );
IBUF  _0733_ (
    .I(m4_data_i[8]),
    .O(_0045_[8])
  );
IBUF  _0734_ (
    .I(m4_data_i[9]),
    .O(_0045_[9])
  );
OBUF  _0735_ (
    .I(_0046_[0]),
    .O(m4_data_o[0])
  );
OBUF  _0736_ (
    .I(_0046_[1]),
    .O(m4_data_o[1])
  );
OBUF  _0737_ (
    .I(_0046_[10]),
    .O(m4_data_o[10])
  );
OBUF  _0738_ (
    .I(_0046_[11]),
    .O(m4_data_o[11])
  );
OBUF  _0739_ (
    .I(_0046_[12]),
    .O(m4_data_o[12])
  );
OBUF  _0740_ (
    .I(_0046_[13]),
    .O(m4_data_o[13])
  );
OBUF  _0741_ (
    .I(_0046_[14]),
    .O(m4_data_o[14])
  );
OBUF  _0742_ (
    .I(_0046_[15]),
    .O(m4_data_o[15])
  );
OBUF  _0743_ (
    .I(_0046_[16]),
    .O(m4_data_o[16])
  );
OBUF  _0744_ (
    .I(_0046_[17]),
    .O(m4_data_o[17])
  );
OBUF  _0745_ (
    .I(_0046_[18]),
    .O(m4_data_o[18])
  );
OBUF  _0746_ (
    .I(_0046_[19]),
    .O(m4_data_o[19])
  );
OBUF  _0747_ (
    .I(_0046_[2]),
    .O(m4_data_o[2])
  );
OBUF  _0748_ (
    .I(_0046_[20]),
    .O(m4_data_o[20])
  );
OBUF  _0749_ (
    .I(_0046_[21]),
    .O(m4_data_o[21])
  );
OBUF  _0750_ (
    .I(_0046_[22]),
    .O(m4_data_o[22])
  );
OBUF  _0751_ (
    .I(_0046_[23]),
    .O(m4_data_o[23])
  );
OBUF  _0752_ (
    .I(_0046_[24]),
    .O(m4_data_o[24])
  );
OBUF  _0753_ (
    .I(_0046_[25]),
    .O(m4_data_o[25])
  );
OBUF  _0754_ (
    .I(_0046_[26]),
    .O(m4_data_o[26])
  );
OBUF  _0755_ (
    .I(_0046_[27]),
    .O(m4_data_o[27])
  );
OBUF  _0756_ (
    .I(_0046_[28]),
    .O(m4_data_o[28])
  );
OBUF  _0757_ (
    .I(_0046_[29]),
    .O(m4_data_o[29])
  );
OBUF  _0758_ (
    .I(_0046_[3]),
    .O(m4_data_o[3])
  );
OBUF  _0759_ (
    .I(_0046_[30]),
    .O(m4_data_o[30])
  );
OBUF  _0760_ (
    .I(_0046_[31]),
    .O(m4_data_o[31])
  );
OBUF  _0761_ (
    .I(_0046_[4]),
    .O(m4_data_o[4])
  );
OBUF  _0762_ (
    .I(_0046_[5]),
    .O(m4_data_o[5])
  );
OBUF  _0763_ (
    .I(_0046_[6]),
    .O(m4_data_o[6])
  );
OBUF  _0764_ (
    .I(_0046_[7]),
    .O(m4_data_o[7])
  );
OBUF  _0765_ (
    .I(_0046_[8]),
    .O(m4_data_o[8])
  );
OBUF  _0766_ (
    .I(_0046_[9]),
    .O(m4_data_o[9])
  );
OBUF  _0767_ (
    .I(_0047_),
    .O(m4_err_o)
  );
OBUF  _0768_ (
    .I(_0048_),
    .O(m4_rty_o)
  );
IBUF  _0769_ (
    .I(m4_sel_i[0]),
    .O(_0049_[0])
  );
IBUF  _0770_ (
    .I(m4_sel_i[1]),
    .O(_0049_[1])
  );
IBUF  _0771_ (
    .I(m4_sel_i[2]),
    .O(_0049_[2])
  );
IBUF  _0772_ (
    .I(m4_sel_i[3]),
    .O(_0049_[3])
  );
IBUF  _0773_ (
    .I(m4_stb_i),
    .O(_0050_)
  );
IBUF  _0774_ (
    .I(m4_we_i),
    .O(_0051_)
  );
OBUF  _0775_ (
    .I(_0052_),
    .O(m5_ack_o)
  );
IBUF  _0776_ (
    .I(m5_addr_i[0]),
    .O(_0053_[0])
  );
IBUF  _0777_ (
    .I(m5_addr_i[1]),
    .O(_0053_[1])
  );
IBUF  _0778_ (
    .I(m5_addr_i[10]),
    .O(_0053_[10])
  );
IBUF  _0779_ (
    .I(m5_addr_i[11]),
    .O(_0053_[11])
  );
IBUF  _0780_ (
    .I(m5_addr_i[12]),
    .O(_0053_[12])
  );
IBUF  _0781_ (
    .I(m5_addr_i[13]),
    .O(_0053_[13])
  );
IBUF  _0782_ (
    .I(m5_addr_i[14]),
    .O(_0053_[14])
  );
IBUF  _0783_ (
    .I(m5_addr_i[15]),
    .O(_0053_[15])
  );
IBUF  _0784_ (
    .I(m5_addr_i[16]),
    .O(_0053_[16])
  );
IBUF  _0785_ (
    .I(m5_addr_i[17]),
    .O(_0053_[17])
  );
IBUF  _0786_ (
    .I(m5_addr_i[18]),
    .O(_0053_[18])
  );
IBUF  _0787_ (
    .I(m5_addr_i[19]),
    .O(_0053_[19])
  );
IBUF  _0788_ (
    .I(m5_addr_i[2]),
    .O(_0053_[2])
  );
IBUF  _0789_ (
    .I(m5_addr_i[20]),
    .O(_0053_[20])
  );
IBUF  _0790_ (
    .I(m5_addr_i[21]),
    .O(_0053_[21])
  );
IBUF  _0791_ (
    .I(m5_addr_i[22]),
    .O(_0053_[22])
  );
IBUF  _0792_ (
    .I(m5_addr_i[23]),
    .O(_0053_[23])
  );
IBUF  _0793_ (
    .I(m5_addr_i[24]),
    .O(_0053_[24])
  );
IBUF  _0794_ (
    .I(m5_addr_i[25]),
    .O(_0053_[25])
  );
IBUF  _0795_ (
    .I(m5_addr_i[26]),
    .O(_0053_[26])
  );
IBUF  _0796_ (
    .I(m5_addr_i[27]),
    .O(_0053_[27])
  );
IBUF  _0797_ (
    .I(m5_addr_i[28]),
    .O(_0053_[28])
  );
IBUF  _0798_ (
    .I(m5_addr_i[29]),
    .O(_0053_[29])
  );
IBUF  _0799_ (
    .I(m5_addr_i[3]),
    .O(_0053_[3])
  );
IBUF  _0800_ (
    .I(m5_addr_i[30]),
    .O(_0053_[30])
  );
IBUF  _0801_ (
    .I(m5_addr_i[31]),
    .O(_0053_[31])
  );
IBUF  _0802_ (
    .I(m5_addr_i[4]),
    .O(_0053_[4])
  );
IBUF  _0803_ (
    .I(m5_addr_i[5]),
    .O(_0053_[5])
  );
IBUF  _0804_ (
    .I(m5_addr_i[6]),
    .O(_0053_[6])
  );
IBUF  _0805_ (
    .I(m5_addr_i[7]),
    .O(_0053_[7])
  );
IBUF  _0806_ (
    .I(m5_addr_i[8]),
    .O(_0053_[8])
  );
IBUF  _0807_ (
    .I(m5_addr_i[9]),
    .O(_0053_[9])
  );
IBUF  _0808_ (
    .I(m5_cyc_i),
    .O(_0054_)
  );
IBUF  _0809_ (
    .I(m5_data_i[0]),
    .O(_0055_[0])
  );
IBUF  _0810_ (
    .I(m5_data_i[1]),
    .O(_0055_[1])
  );
IBUF  _0811_ (
    .I(m5_data_i[10]),
    .O(_0055_[10])
  );
IBUF  _0812_ (
    .I(m5_data_i[11]),
    .O(_0055_[11])
  );
IBUF  _0813_ (
    .I(m5_data_i[12]),
    .O(_0055_[12])
  );
IBUF  _0814_ (
    .I(m5_data_i[13]),
    .O(_0055_[13])
  );
IBUF  _0815_ (
    .I(m5_data_i[14]),
    .O(_0055_[14])
  );
IBUF  _0816_ (
    .I(m5_data_i[15]),
    .O(_0055_[15])
  );
IBUF  _0817_ (
    .I(m5_data_i[16]),
    .O(_0055_[16])
  );
IBUF  _0818_ (
    .I(m5_data_i[17]),
    .O(_0055_[17])
  );
IBUF  _0819_ (
    .I(m5_data_i[18]),
    .O(_0055_[18])
  );
IBUF  _0820_ (
    .I(m5_data_i[19]),
    .O(_0055_[19])
  );
IBUF  _0821_ (
    .I(m5_data_i[2]),
    .O(_0055_[2])
  );
IBUF  _0822_ (
    .I(m5_data_i[20]),
    .O(_0055_[20])
  );
IBUF  _0823_ (
    .I(m5_data_i[21]),
    .O(_0055_[21])
  );
IBUF  _0824_ (
    .I(m5_data_i[22]),
    .O(_0055_[22])
  );
IBUF  _0825_ (
    .I(m5_data_i[23]),
    .O(_0055_[23])
  );
IBUF  _0826_ (
    .I(m5_data_i[24]),
    .O(_0055_[24])
  );
IBUF  _0827_ (
    .I(m5_data_i[25]),
    .O(_0055_[25])
  );
IBUF  _0828_ (
    .I(m5_data_i[26]),
    .O(_0055_[26])
  );
IBUF  _0829_ (
    .I(m5_data_i[27]),
    .O(_0055_[27])
  );
IBUF  _0830_ (
    .I(m5_data_i[28]),
    .O(_0055_[28])
  );
IBUF  _0831_ (
    .I(m5_data_i[29]),
    .O(_0055_[29])
  );
IBUF  _0832_ (
    .I(m5_data_i[3]),
    .O(_0055_[3])
  );
IBUF  _0833_ (
    .I(m5_data_i[30]),
    .O(_0055_[30])
  );
IBUF  _0834_ (
    .I(m5_data_i[31]),
    .O(_0055_[31])
  );
IBUF  _0835_ (
    .I(m5_data_i[4]),
    .O(_0055_[4])
  );
IBUF  _0836_ (
    .I(m5_data_i[5]),
    .O(_0055_[5])
  );
IBUF  _0837_ (
    .I(m5_data_i[6]),
    .O(_0055_[6])
  );
IBUF  _0838_ (
    .I(m5_data_i[7]),
    .O(_0055_[7])
  );
IBUF  _0839_ (
    .I(m5_data_i[8]),
    .O(_0055_[8])
  );
IBUF  _0840_ (
    .I(m5_data_i[9]),
    .O(_0055_[9])
  );
OBUF  _0841_ (
    .I(_0056_[0]),
    .O(m5_data_o[0])
  );
OBUF  _0842_ (
    .I(_0056_[1]),
    .O(m5_data_o[1])
  );
OBUF  _0843_ (
    .I(_0056_[10]),
    .O(m5_data_o[10])
  );
OBUF  _0844_ (
    .I(_0056_[11]),
    .O(m5_data_o[11])
  );
OBUF  _0845_ (
    .I(_0056_[12]),
    .O(m5_data_o[12])
  );
OBUF  _0846_ (
    .I(_0056_[13]),
    .O(m5_data_o[13])
  );
OBUF  _0847_ (
    .I(_0056_[14]),
    .O(m5_data_o[14])
  );
OBUF  _0848_ (
    .I(_0056_[15]),
    .O(m5_data_o[15])
  );
OBUF  _0849_ (
    .I(_0056_[16]),
    .O(m5_data_o[16])
  );
OBUF  _0850_ (
    .I(_0056_[17]),
    .O(m5_data_o[17])
  );
OBUF  _0851_ (
    .I(_0056_[18]),
    .O(m5_data_o[18])
  );
OBUF  _0852_ (
    .I(_0056_[19]),
    .O(m5_data_o[19])
  );
OBUF  _0853_ (
    .I(_0056_[2]),
    .O(m5_data_o[2])
  );
OBUF  _0854_ (
    .I(_0056_[20]),
    .O(m5_data_o[20])
  );
OBUF  _0855_ (
    .I(_0056_[21]),
    .O(m5_data_o[21])
  );
OBUF  _0856_ (
    .I(_0056_[22]),
    .O(m5_data_o[22])
  );
OBUF  _0857_ (
    .I(_0056_[23]),
    .O(m5_data_o[23])
  );
OBUF  _0858_ (
    .I(_0056_[24]),
    .O(m5_data_o[24])
  );
OBUF  _0859_ (
    .I(_0056_[25]),
    .O(m5_data_o[25])
  );
OBUF  _0860_ (
    .I(_0056_[26]),
    .O(m5_data_o[26])
  );
OBUF  _0861_ (
    .I(_0056_[27]),
    .O(m5_data_o[27])
  );
OBUF  _0862_ (
    .I(_0056_[28]),
    .O(m5_data_o[28])
  );
OBUF  _0863_ (
    .I(_0056_[29]),
    .O(m5_data_o[29])
  );
OBUF  _0864_ (
    .I(_0056_[3]),
    .O(m5_data_o[3])
  );
OBUF  _0865_ (
    .I(_0056_[30]),
    .O(m5_data_o[30])
  );
OBUF  _0866_ (
    .I(_0056_[31]),
    .O(m5_data_o[31])
  );
OBUF  _0867_ (
    .I(_0056_[4]),
    .O(m5_data_o[4])
  );
OBUF  _0868_ (
    .I(_0056_[5]),
    .O(m5_data_o[5])
  );
OBUF  _0869_ (
    .I(_0056_[6]),
    .O(m5_data_o[6])
  );
OBUF  _0870_ (
    .I(_0056_[7]),
    .O(m5_data_o[7])
  );
OBUF  _0871_ (
    .I(_0056_[8]),
    .O(m5_data_o[8])
  );
OBUF  _0872_ (
    .I(_0056_[9]),
    .O(m5_data_o[9])
  );
OBUF  _0873_ (
    .I(_0057_),
    .O(m5_err_o)
  );
OBUF  _0874_ (
    .I(_0058_),
    .O(m5_rty_o)
  );
IBUF  _0875_ (
    .I(m5_sel_i[0]),
    .O(_0059_[0])
  );
IBUF  _0876_ (
    .I(m5_sel_i[1]),
    .O(_0059_[1])
  );
IBUF  _0877_ (
    .I(m5_sel_i[2]),
    .O(_0059_[2])
  );
IBUF  _0878_ (
    .I(m5_sel_i[3]),
    .O(_0059_[3])
  );
IBUF  _0879_ (
    .I(m5_stb_i),
    .O(_0060_)
  );
IBUF  _0880_ (
    .I(m5_we_i),
    .O(_0061_)
  );
OBUF  _0881_ (
    .I(_0062_),
    .O(m6_ack_o)
  );
IBUF  _0882_ (
    .I(m6_addr_i[0]),
    .O(_0063_[0])
  );
IBUF  _0883_ (
    .I(m6_addr_i[1]),
    .O(_0063_[1])
  );
IBUF  _0884_ (
    .I(m6_addr_i[10]),
    .O(_0063_[10])
  );
IBUF  _0885_ (
    .I(m6_addr_i[11]),
    .O(_0063_[11])
  );
IBUF  _0886_ (
    .I(m6_addr_i[12]),
    .O(_0063_[12])
  );
IBUF  _0887_ (
    .I(m6_addr_i[13]),
    .O(_0063_[13])
  );
IBUF  _0888_ (
    .I(m6_addr_i[14]),
    .O(_0063_[14])
  );
IBUF  _0889_ (
    .I(m6_addr_i[15]),
    .O(_0063_[15])
  );
IBUF  _0890_ (
    .I(m6_addr_i[16]),
    .O(_0063_[16])
  );
IBUF  _0891_ (
    .I(m6_addr_i[17]),
    .O(_0063_[17])
  );
IBUF  _0892_ (
    .I(m6_addr_i[18]),
    .O(_0063_[18])
  );
IBUF  _0893_ (
    .I(m6_addr_i[19]),
    .O(_0063_[19])
  );
IBUF  _0894_ (
    .I(m6_addr_i[2]),
    .O(_0063_[2])
  );
IBUF  _0895_ (
    .I(m6_addr_i[20]),
    .O(_0063_[20])
  );
IBUF  _0896_ (
    .I(m6_addr_i[21]),
    .O(_0063_[21])
  );
IBUF  _0897_ (
    .I(m6_addr_i[22]),
    .O(_0063_[22])
  );
IBUF  _0898_ (
    .I(m6_addr_i[23]),
    .O(_0063_[23])
  );
IBUF  _0899_ (
    .I(m6_addr_i[24]),
    .O(_0063_[24])
  );
IBUF  _0900_ (
    .I(m6_addr_i[25]),
    .O(_0063_[25])
  );
IBUF  _0901_ (
    .I(m6_addr_i[26]),
    .O(_0063_[26])
  );
IBUF  _0902_ (
    .I(m6_addr_i[27]),
    .O(_0063_[27])
  );
IBUF  _0903_ (
    .I(m6_addr_i[28]),
    .O(_0063_[28])
  );
IBUF  _0904_ (
    .I(m6_addr_i[29]),
    .O(_0063_[29])
  );
IBUF  _0905_ (
    .I(m6_addr_i[3]),
    .O(_0063_[3])
  );
IBUF  _0906_ (
    .I(m6_addr_i[30]),
    .O(_0063_[30])
  );
IBUF  _0907_ (
    .I(m6_addr_i[31]),
    .O(_0063_[31])
  );
IBUF  _0908_ (
    .I(m6_addr_i[4]),
    .O(_0063_[4])
  );
IBUF  _0909_ (
    .I(m6_addr_i[5]),
    .O(_0063_[5])
  );
IBUF  _0910_ (
    .I(m6_addr_i[6]),
    .O(_0063_[6])
  );
IBUF  _0911_ (
    .I(m6_addr_i[7]),
    .O(_0063_[7])
  );
IBUF  _0912_ (
    .I(m6_addr_i[8]),
    .O(_0063_[8])
  );
IBUF  _0913_ (
    .I(m6_addr_i[9]),
    .O(_0063_[9])
  );
IBUF  _0914_ (
    .I(m6_cyc_i),
    .O(_0064_)
  );
IBUF  _0915_ (
    .I(m6_data_i[0]),
    .O(_0065_[0])
  );
IBUF  _0916_ (
    .I(m6_data_i[1]),
    .O(_0065_[1])
  );
IBUF  _0917_ (
    .I(m6_data_i[10]),
    .O(_0065_[10])
  );
IBUF  _0918_ (
    .I(m6_data_i[11]),
    .O(_0065_[11])
  );
IBUF  _0919_ (
    .I(m6_data_i[12]),
    .O(_0065_[12])
  );
IBUF  _0920_ (
    .I(m6_data_i[13]),
    .O(_0065_[13])
  );
IBUF  _0921_ (
    .I(m6_data_i[14]),
    .O(_0065_[14])
  );
IBUF  _0922_ (
    .I(m6_data_i[15]),
    .O(_0065_[15])
  );
IBUF  _0923_ (
    .I(m6_data_i[16]),
    .O(_0065_[16])
  );
IBUF  _0924_ (
    .I(m6_data_i[17]),
    .O(_0065_[17])
  );
IBUF  _0925_ (
    .I(m6_data_i[18]),
    .O(_0065_[18])
  );
IBUF  _0926_ (
    .I(m6_data_i[19]),
    .O(_0065_[19])
  );
IBUF  _0927_ (
    .I(m6_data_i[2]),
    .O(_0065_[2])
  );
IBUF  _0928_ (
    .I(m6_data_i[20]),
    .O(_0065_[20])
  );
IBUF  _0929_ (
    .I(m6_data_i[21]),
    .O(_0065_[21])
  );
IBUF  _0930_ (
    .I(m6_data_i[22]),
    .O(_0065_[22])
  );
IBUF  _0931_ (
    .I(m6_data_i[23]),
    .O(_0065_[23])
  );
IBUF  _0932_ (
    .I(m6_data_i[24]),
    .O(_0065_[24])
  );
IBUF  _0933_ (
    .I(m6_data_i[25]),
    .O(_0065_[25])
  );
IBUF  _0934_ (
    .I(m6_data_i[26]),
    .O(_0065_[26])
  );
IBUF  _0935_ (
    .I(m6_data_i[27]),
    .O(_0065_[27])
  );
IBUF  _0936_ (
    .I(m6_data_i[28]),
    .O(_0065_[28])
  );
IBUF  _0937_ (
    .I(m6_data_i[29]),
    .O(_0065_[29])
  );
IBUF  _0938_ (
    .I(m6_data_i[3]),
    .O(_0065_[3])
  );
IBUF  _0939_ (
    .I(m6_data_i[30]),
    .O(_0065_[30])
  );
IBUF  _0940_ (
    .I(m6_data_i[31]),
    .O(_0065_[31])
  );
IBUF  _0941_ (
    .I(m6_data_i[4]),
    .O(_0065_[4])
  );
IBUF  _0942_ (
    .I(m6_data_i[5]),
    .O(_0065_[5])
  );
IBUF  _0943_ (
    .I(m6_data_i[6]),
    .O(_0065_[6])
  );
IBUF  _0944_ (
    .I(m6_data_i[7]),
    .O(_0065_[7])
  );
IBUF  _0945_ (
    .I(m6_data_i[8]),
    .O(_0065_[8])
  );
IBUF  _0946_ (
    .I(m6_data_i[9]),
    .O(_0065_[9])
  );
OBUF  _0947_ (
    .I(_0066_[0]),
    .O(m6_data_o[0])
  );
OBUF  _0948_ (
    .I(_0066_[1]),
    .O(m6_data_o[1])
  );
OBUF  _0949_ (
    .I(_0066_[10]),
    .O(m6_data_o[10])
  );
OBUF  _0950_ (
    .I(_0066_[11]),
    .O(m6_data_o[11])
  );
OBUF  _0951_ (
    .I(_0066_[12]),
    .O(m6_data_o[12])
  );
OBUF  _0952_ (
    .I(_0066_[13]),
    .O(m6_data_o[13])
  );
OBUF  _0953_ (
    .I(_0066_[14]),
    .O(m6_data_o[14])
  );
OBUF  _0954_ (
    .I(_0066_[15]),
    .O(m6_data_o[15])
  );
OBUF  _0955_ (
    .I(_0066_[16]),
    .O(m6_data_o[16])
  );
OBUF  _0956_ (
    .I(_0066_[17]),
    .O(m6_data_o[17])
  );
OBUF  _0957_ (
    .I(_0066_[18]),
    .O(m6_data_o[18])
  );
OBUF  _0958_ (
    .I(_0066_[19]),
    .O(m6_data_o[19])
  );
OBUF  _0959_ (
    .I(_0066_[2]),
    .O(m6_data_o[2])
  );
OBUF  _0960_ (
    .I(_0066_[20]),
    .O(m6_data_o[20])
  );
OBUF  _0961_ (
    .I(_0066_[21]),
    .O(m6_data_o[21])
  );
OBUF  _0962_ (
    .I(_0066_[22]),
    .O(m6_data_o[22])
  );
OBUF  _0963_ (
    .I(_0066_[23]),
    .O(m6_data_o[23])
  );
OBUF  _0964_ (
    .I(_0066_[24]),
    .O(m6_data_o[24])
  );
OBUF  _0965_ (
    .I(_0066_[25]),
    .O(m6_data_o[25])
  );
OBUF  _0966_ (
    .I(_0066_[26]),
    .O(m6_data_o[26])
  );
OBUF  _0967_ (
    .I(_0066_[27]),
    .O(m6_data_o[27])
  );
OBUF  _0968_ (
    .I(_0066_[28]),
    .O(m6_data_o[28])
  );
OBUF  _0969_ (
    .I(_0066_[29]),
    .O(m6_data_o[29])
  );
OBUF  _0970_ (
    .I(_0066_[3]),
    .O(m6_data_o[3])
  );
OBUF  _0971_ (
    .I(_0066_[30]),
    .O(m6_data_o[30])
  );
OBUF  _0972_ (
    .I(_0066_[31]),
    .O(m6_data_o[31])
  );
OBUF  _0973_ (
    .I(_0066_[4]),
    .O(m6_data_o[4])
  );
OBUF  _0974_ (
    .I(_0066_[5]),
    .O(m6_data_o[5])
  );
OBUF  _0975_ (
    .I(_0066_[6]),
    .O(m6_data_o[6])
  );
OBUF  _0976_ (
    .I(_0066_[7]),
    .O(m6_data_o[7])
  );
OBUF  _0977_ (
    .I(_0066_[8]),
    .O(m6_data_o[8])
  );
OBUF  _0978_ (
    .I(_0066_[9]),
    .O(m6_data_o[9])
  );
OBUF  _0979_ (
    .I(_0067_),
    .O(m6_err_o)
  );
OBUF  _0980_ (
    .I(_0068_),
    .O(m6_rty_o)
  );
IBUF  _0981_ (
    .I(m6_sel_i[0]),
    .O(_0069_[0])
  );
IBUF  _0982_ (
    .I(m6_sel_i[1]),
    .O(_0069_[1])
  );
IBUF  _0983_ (
    .I(m6_sel_i[2]),
    .O(_0069_[2])
  );
IBUF  _0984_ (
    .I(m6_sel_i[3]),
    .O(_0069_[3])
  );
IBUF  _0985_ (
    .I(m6_stb_i),
    .O(_0070_)
  );
IBUF  _0986_ (
    .I(m6_we_i),
    .O(_0071_)
  );
OBUF  _0987_ (
    .I(_0072_),
    .O(m7_ack_o)
  );
IBUF  _0988_ (
    .I(m7_addr_i[0]),
    .O(_0073_[0])
  );
IBUF  _0989_ (
    .I(m7_addr_i[1]),
    .O(_0073_[1])
  );
IBUF  _0990_ (
    .I(m7_addr_i[10]),
    .O(_0073_[10])
  );
IBUF  _0991_ (
    .I(m7_addr_i[11]),
    .O(_0073_[11])
  );
IBUF  _0992_ (
    .I(m7_addr_i[12]),
    .O(_0073_[12])
  );
IBUF  _0993_ (
    .I(m7_addr_i[13]),
    .O(_0073_[13])
  );
IBUF  _0994_ (
    .I(m7_addr_i[14]),
    .O(_0073_[14])
  );
IBUF  _0995_ (
    .I(m7_addr_i[15]),
    .O(_0073_[15])
  );
IBUF  _0996_ (
    .I(m7_addr_i[16]),
    .O(_0073_[16])
  );
IBUF  _0997_ (
    .I(m7_addr_i[17]),
    .O(_0073_[17])
  );
IBUF  _0998_ (
    .I(m7_addr_i[18]),
    .O(_0073_[18])
  );
IBUF  _0999_ (
    .I(m7_addr_i[19]),
    .O(_0073_[19])
  );
IBUF  _1000_ (
    .I(m7_addr_i[2]),
    .O(_0073_[2])
  );
IBUF  _1001_ (
    .I(m7_addr_i[20]),
    .O(_0073_[20])
  );
IBUF  _1002_ (
    .I(m7_addr_i[21]),
    .O(_0073_[21])
  );
IBUF  _1003_ (
    .I(m7_addr_i[22]),
    .O(_0073_[22])
  );
IBUF  _1004_ (
    .I(m7_addr_i[23]),
    .O(_0073_[23])
  );
IBUF  _1005_ (
    .I(m7_addr_i[24]),
    .O(_0073_[24])
  );
IBUF  _1006_ (
    .I(m7_addr_i[25]),
    .O(_0073_[25])
  );
IBUF  _1007_ (
    .I(m7_addr_i[26]),
    .O(_0073_[26])
  );
IBUF  _1008_ (
    .I(m7_addr_i[27]),
    .O(_0073_[27])
  );
IBUF  _1009_ (
    .I(m7_addr_i[28]),
    .O(_0073_[28])
  );
IBUF  _1010_ (
    .I(m7_addr_i[29]),
    .O(_0073_[29])
  );
IBUF  _1011_ (
    .I(m7_addr_i[3]),
    .O(_0073_[3])
  );
IBUF  _1012_ (
    .I(m7_addr_i[30]),
    .O(_0073_[30])
  );
IBUF  _1013_ (
    .I(m7_addr_i[31]),
    .O(_0073_[31])
  );
IBUF  _1014_ (
    .I(m7_addr_i[4]),
    .O(_0073_[4])
  );
IBUF  _1015_ (
    .I(m7_addr_i[5]),
    .O(_0073_[5])
  );
IBUF  _1016_ (
    .I(m7_addr_i[6]),
    .O(_0073_[6])
  );
IBUF  _1017_ (
    .I(m7_addr_i[7]),
    .O(_0073_[7])
  );
IBUF  _1018_ (
    .I(m7_addr_i[8]),
    .O(_0073_[8])
  );
IBUF  _1019_ (
    .I(m7_addr_i[9]),
    .O(_0073_[9])
  );
IBUF  _1020_ (
    .I(m7_cyc_i),
    .O(_0074_)
  );
IBUF  _1021_ (
    .I(m7_data_i[0]),
    .O(_0075_[0])
  );
IBUF  _1022_ (
    .I(m7_data_i[1]),
    .O(_0075_[1])
  );
IBUF  _1023_ (
    .I(m7_data_i[10]),
    .O(_0075_[10])
  );
IBUF  _1024_ (
    .I(m7_data_i[11]),
    .O(_0075_[11])
  );
IBUF  _1025_ (
    .I(m7_data_i[12]),
    .O(_0075_[12])
  );
IBUF  _1026_ (
    .I(m7_data_i[13]),
    .O(_0075_[13])
  );
IBUF  _1027_ (
    .I(m7_data_i[14]),
    .O(_0075_[14])
  );
IBUF  _1028_ (
    .I(m7_data_i[15]),
    .O(_0075_[15])
  );
IBUF  _1029_ (
    .I(m7_data_i[16]),
    .O(_0075_[16])
  );
IBUF  _1030_ (
    .I(m7_data_i[17]),
    .O(_0075_[17])
  );
IBUF  _1031_ (
    .I(m7_data_i[18]),
    .O(_0075_[18])
  );
IBUF  _1032_ (
    .I(m7_data_i[19]),
    .O(_0075_[19])
  );
IBUF  _1033_ (
    .I(m7_data_i[2]),
    .O(_0075_[2])
  );
IBUF  _1034_ (
    .I(m7_data_i[20]),
    .O(_0075_[20])
  );
IBUF  _1035_ (
    .I(m7_data_i[21]),
    .O(_0075_[21])
  );
IBUF  _1036_ (
    .I(m7_data_i[22]),
    .O(_0075_[22])
  );
IBUF  _1037_ (
    .I(m7_data_i[23]),
    .O(_0075_[23])
  );
IBUF  _1038_ (
    .I(m7_data_i[24]),
    .O(_0075_[24])
  );
IBUF  _1039_ (
    .I(m7_data_i[25]),
    .O(_0075_[25])
  );
IBUF  _1040_ (
    .I(m7_data_i[26]),
    .O(_0075_[26])
  );
IBUF  _1041_ (
    .I(m7_data_i[27]),
    .O(_0075_[27])
  );
IBUF  _1042_ (
    .I(m7_data_i[28]),
    .O(_0075_[28])
  );
IBUF  _1043_ (
    .I(m7_data_i[29]),
    .O(_0075_[29])
  );
IBUF  _1044_ (
    .I(m7_data_i[3]),
    .O(_0075_[3])
  );
IBUF  _1045_ (
    .I(m7_data_i[30]),
    .O(_0075_[30])
  );
IBUF  _1046_ (
    .I(m7_data_i[31]),
    .O(_0075_[31])
  );
IBUF  _1047_ (
    .I(m7_data_i[4]),
    .O(_0075_[4])
  );
IBUF  _1048_ (
    .I(m7_data_i[5]),
    .O(_0075_[5])
  );
IBUF  _1049_ (
    .I(m7_data_i[6]),
    .O(_0075_[6])
  );
IBUF  _1050_ (
    .I(m7_data_i[7]),
    .O(_0075_[7])
  );
IBUF  _1051_ (
    .I(m7_data_i[8]),
    .O(_0075_[8])
  );
IBUF  _1052_ (
    .I(m7_data_i[9]),
    .O(_0075_[9])
  );
OBUF  _1053_ (
    .I(_0076_[0]),
    .O(m7_data_o[0])
  );
OBUF  _1054_ (
    .I(_0076_[1]),
    .O(m7_data_o[1])
  );
OBUF  _1055_ (
    .I(_0076_[10]),
    .O(m7_data_o[10])
  );
OBUF  _1056_ (
    .I(_0076_[11]),
    .O(m7_data_o[11])
  );
OBUF  _1057_ (
    .I(_0076_[12]),
    .O(m7_data_o[12])
  );
OBUF  _1058_ (
    .I(_0076_[13]),
    .O(m7_data_o[13])
  );
OBUF  _1059_ (
    .I(_0076_[14]),
    .O(m7_data_o[14])
  );
OBUF  _1060_ (
    .I(_0076_[15]),
    .O(m7_data_o[15])
  );
OBUF  _1061_ (
    .I(_0076_[16]),
    .O(m7_data_o[16])
  );
OBUF  _1062_ (
    .I(_0076_[17]),
    .O(m7_data_o[17])
  );
OBUF  _1063_ (
    .I(_0076_[18]),
    .O(m7_data_o[18])
  );
OBUF  _1064_ (
    .I(_0076_[19]),
    .O(m7_data_o[19])
  );
OBUF  _1065_ (
    .I(_0076_[2]),
    .O(m7_data_o[2])
  );
OBUF  _1066_ (
    .I(_0076_[20]),
    .O(m7_data_o[20])
  );
OBUF  _1067_ (
    .I(_0076_[21]),
    .O(m7_data_o[21])
  );
OBUF  _1068_ (
    .I(_0076_[22]),
    .O(m7_data_o[22])
  );
OBUF  _1069_ (
    .I(_0076_[23]),
    .O(m7_data_o[23])
  );
OBUF  _1070_ (
    .I(_0076_[24]),
    .O(m7_data_o[24])
  );
OBUF  _1071_ (
    .I(_0076_[25]),
    .O(m7_data_o[25])
  );
OBUF  _1072_ (
    .I(_0076_[26]),
    .O(m7_data_o[26])
  );
OBUF  _1073_ (
    .I(_0076_[27]),
    .O(m7_data_o[27])
  );
OBUF  _1074_ (
    .I(_0076_[28]),
    .O(m7_data_o[28])
  );
OBUF  _1075_ (
    .I(_0076_[29]),
    .O(m7_data_o[29])
  );
OBUF  _1076_ (
    .I(_0076_[3]),
    .O(m7_data_o[3])
  );
OBUF  _1077_ (
    .I(_0076_[30]),
    .O(m7_data_o[30])
  );
OBUF  _1078_ (
    .I(_0076_[31]),
    .O(m7_data_o[31])
  );
OBUF  _1079_ (
    .I(_0076_[4]),
    .O(m7_data_o[4])
  );
OBUF  _1080_ (
    .I(_0076_[5]),
    .O(m7_data_o[5])
  );
OBUF  _1081_ (
    .I(_0076_[6]),
    .O(m7_data_o[6])
  );
OBUF  _1082_ (
    .I(_0076_[7]),
    .O(m7_data_o[7])
  );
OBUF  _1083_ (
    .I(_0076_[8]),
    .O(m7_data_o[8])
  );
OBUF  _1084_ (
    .I(_0076_[9]),
    .O(m7_data_o[9])
  );
OBUF  _1085_ (
    .I(_0077_),
    .O(m7_err_o)
  );
OBUF  _1086_ (
    .I(_0078_),
    .O(m7_rty_o)
  );
IBUF  _1087_ (
    .I(m7_sel_i[0]),
    .O(_0079_[0])
  );
IBUF  _1088_ (
    .I(m7_sel_i[1]),
    .O(_0079_[1])
  );
IBUF  _1089_ (
    .I(m7_sel_i[2]),
    .O(_0079_[2])
  );
IBUF  _1090_ (
    .I(m7_sel_i[3]),
    .O(_0079_[3])
  );
IBUF  _1091_ (
    .I(m7_stb_i),
    .O(_0080_)
  );
IBUF  _1092_ (
    .I(m7_we_i),
    .O(_0081_)
  );
IBUF  _1093_ (
    .I(rst_i),
    .O(_0082_)
  );
IBUF  _1094_ (
    .I(s0_ack_i),
    .O(_0083_)
  );
OBUF  _1095_ (
    .I(_0084_[0]),
    .O(s0_addr_o[0])
  );
OBUF  _1096_ (
    .I(_0084_[1]),
    .O(s0_addr_o[1])
  );
OBUF  _1097_ (
    .I(_0084_[10]),
    .O(s0_addr_o[10])
  );
OBUF  _1098_ (
    .I(_0084_[11]),
    .O(s0_addr_o[11])
  );
OBUF  _1099_ (
    .I(_0084_[12]),
    .O(s0_addr_o[12])
  );
OBUF  _1100_ (
    .I(_0084_[13]),
    .O(s0_addr_o[13])
  );
OBUF  _1101_ (
    .I(_0084_[14]),
    .O(s0_addr_o[14])
  );
OBUF  _1102_ (
    .I(_0084_[15]),
    .O(s0_addr_o[15])
  );
OBUF  _1103_ (
    .I(_0084_[16]),
    .O(s0_addr_o[16])
  );
OBUF  _1104_ (
    .I(_0084_[17]),
    .O(s0_addr_o[17])
  );
OBUF  _1105_ (
    .I(_0084_[18]),
    .O(s0_addr_o[18])
  );
OBUF  _1106_ (
    .I(_0084_[19]),
    .O(s0_addr_o[19])
  );
OBUF  _1107_ (
    .I(_0084_[2]),
    .O(s0_addr_o[2])
  );
OBUF  _1108_ (
    .I(_0084_[20]),
    .O(s0_addr_o[20])
  );
OBUF  _1109_ (
    .I(_0084_[21]),
    .O(s0_addr_o[21])
  );
OBUF  _1110_ (
    .I(_0084_[22]),
    .O(s0_addr_o[22])
  );
OBUF  _1111_ (
    .I(_0084_[23]),
    .O(s0_addr_o[23])
  );
OBUF  _1112_ (
    .I(_0084_[24]),
    .O(s0_addr_o[24])
  );
OBUF  _1113_ (
    .I(_0084_[25]),
    .O(s0_addr_o[25])
  );
OBUF  _1114_ (
    .I(_0084_[26]),
    .O(s0_addr_o[26])
  );
OBUF  _1115_ (
    .I(_0084_[27]),
    .O(s0_addr_o[27])
  );
OBUF  _1116_ (
    .I(_0084_[28]),
    .O(s0_addr_o[28])
  );
OBUF  _1117_ (
    .I(_0084_[29]),
    .O(s0_addr_o[29])
  );
OBUF  _1118_ (
    .I(_0084_[3]),
    .O(s0_addr_o[3])
  );
OBUF  _1119_ (
    .I(_0084_[30]),
    .O(s0_addr_o[30])
  );
OBUF  _1120_ (
    .I(_0084_[31]),
    .O(s0_addr_o[31])
  );
OBUF  _1121_ (
    .I(_0084_[4]),
    .O(s0_addr_o[4])
  );
OBUF  _1122_ (
    .I(_0084_[5]),
    .O(s0_addr_o[5])
  );
OBUF  _1123_ (
    .I(_0084_[6]),
    .O(s0_addr_o[6])
  );
OBUF  _1124_ (
    .I(_0084_[7]),
    .O(s0_addr_o[7])
  );
OBUF  _1125_ (
    .I(_0084_[8]),
    .O(s0_addr_o[8])
  );
OBUF  _1126_ (
    .I(_0084_[9]),
    .O(s0_addr_o[9])
  );
OBUF  _1127_ (
    .I(_0085_),
    .O(s0_cyc_o)
  );
IBUF  _1128_ (
    .I(s0_data_i[0]),
    .O(_0086_[0])
  );
IBUF  _1129_ (
    .I(s0_data_i[1]),
    .O(_0086_[1])
  );
IBUF  _1130_ (
    .I(s0_data_i[10]),
    .O(_0086_[10])
  );
IBUF  _1131_ (
    .I(s0_data_i[11]),
    .O(_0086_[11])
  );
IBUF  _1132_ (
    .I(s0_data_i[12]),
    .O(_0086_[12])
  );
IBUF  _1133_ (
    .I(s0_data_i[13]),
    .O(_0086_[13])
  );
IBUF  _1134_ (
    .I(s0_data_i[14]),
    .O(_0086_[14])
  );
IBUF  _1135_ (
    .I(s0_data_i[15]),
    .O(_0086_[15])
  );
IBUF  _1136_ (
    .I(s0_data_i[16]),
    .O(_0086_[16])
  );
IBUF  _1137_ (
    .I(s0_data_i[17]),
    .O(_0086_[17])
  );
IBUF  _1138_ (
    .I(s0_data_i[18]),
    .O(_0086_[18])
  );
IBUF  _1139_ (
    .I(s0_data_i[19]),
    .O(_0086_[19])
  );
IBUF  _1140_ (
    .I(s0_data_i[2]),
    .O(_0086_[2])
  );
IBUF  _1141_ (
    .I(s0_data_i[20]),
    .O(_0086_[20])
  );
IBUF  _1142_ (
    .I(s0_data_i[21]),
    .O(_0086_[21])
  );
IBUF  _1143_ (
    .I(s0_data_i[22]),
    .O(_0086_[22])
  );
IBUF  _1144_ (
    .I(s0_data_i[23]),
    .O(_0086_[23])
  );
IBUF  _1145_ (
    .I(s0_data_i[24]),
    .O(_0086_[24])
  );
IBUF  _1146_ (
    .I(s0_data_i[25]),
    .O(_0086_[25])
  );
IBUF  _1147_ (
    .I(s0_data_i[26]),
    .O(_0086_[26])
  );
IBUF  _1148_ (
    .I(s0_data_i[27]),
    .O(_0086_[27])
  );
IBUF  _1149_ (
    .I(s0_data_i[28]),
    .O(_0086_[28])
  );
IBUF  _1150_ (
    .I(s0_data_i[29]),
    .O(_0086_[29])
  );
IBUF  _1151_ (
    .I(s0_data_i[3]),
    .O(_0086_[3])
  );
IBUF  _1152_ (
    .I(s0_data_i[30]),
    .O(_0086_[30])
  );
IBUF  _1153_ (
    .I(s0_data_i[31]),
    .O(_0086_[31])
  );
IBUF  _1154_ (
    .I(s0_data_i[4]),
    .O(_0086_[4])
  );
IBUF  _1155_ (
    .I(s0_data_i[5]),
    .O(_0086_[5])
  );
IBUF  _1156_ (
    .I(s0_data_i[6]),
    .O(_0086_[6])
  );
IBUF  _1157_ (
    .I(s0_data_i[7]),
    .O(_0086_[7])
  );
IBUF  _1158_ (
    .I(s0_data_i[8]),
    .O(_0086_[8])
  );
IBUF  _1159_ (
    .I(s0_data_i[9]),
    .O(_0086_[9])
  );
OBUF  _1160_ (
    .I(_0087_[0]),
    .O(s0_data_o[0])
  );
OBUF  _1161_ (
    .I(_0087_[1]),
    .O(s0_data_o[1])
  );
OBUF  _1162_ (
    .I(_0087_[10]),
    .O(s0_data_o[10])
  );
OBUF  _1163_ (
    .I(_0087_[11]),
    .O(s0_data_o[11])
  );
OBUF  _1164_ (
    .I(_0087_[12]),
    .O(s0_data_o[12])
  );
OBUF  _1165_ (
    .I(_0087_[13]),
    .O(s0_data_o[13])
  );
OBUF  _1166_ (
    .I(_0087_[14]),
    .O(s0_data_o[14])
  );
OBUF  _1167_ (
    .I(_0087_[15]),
    .O(s0_data_o[15])
  );
OBUF  _1168_ (
    .I(_0087_[16]),
    .O(s0_data_o[16])
  );
OBUF  _1169_ (
    .I(_0087_[17]),
    .O(s0_data_o[17])
  );
OBUF  _1170_ (
    .I(_0087_[18]),
    .O(s0_data_o[18])
  );
OBUF  _1171_ (
    .I(_0087_[19]),
    .O(s0_data_o[19])
  );
OBUF  _1172_ (
    .I(_0087_[2]),
    .O(s0_data_o[2])
  );
OBUF  _1173_ (
    .I(_0087_[20]),
    .O(s0_data_o[20])
  );
OBUF  _1174_ (
    .I(_0087_[21]),
    .O(s0_data_o[21])
  );
OBUF  _1175_ (
    .I(_0087_[22]),
    .O(s0_data_o[22])
  );
OBUF  _1176_ (
    .I(_0087_[23]),
    .O(s0_data_o[23])
  );
OBUF  _1177_ (
    .I(_0087_[24]),
    .O(s0_data_o[24])
  );
OBUF  _1178_ (
    .I(_0087_[25]),
    .O(s0_data_o[25])
  );
OBUF  _1179_ (
    .I(_0087_[26]),
    .O(s0_data_o[26])
  );
OBUF  _1180_ (
    .I(_0087_[27]),
    .O(s0_data_o[27])
  );
OBUF  _1181_ (
    .I(_0087_[28]),
    .O(s0_data_o[28])
  );
OBUF  _1182_ (
    .I(_0087_[29]),
    .O(s0_data_o[29])
  );
OBUF  _1183_ (
    .I(_0087_[3]),
    .O(s0_data_o[3])
  );
OBUF  _1184_ (
    .I(_0087_[30]),
    .O(s0_data_o[30])
  );
OBUF  _1185_ (
    .I(_0087_[31]),
    .O(s0_data_o[31])
  );
OBUF  _1186_ (
    .I(_0087_[4]),
    .O(s0_data_o[4])
  );
OBUF  _1187_ (
    .I(_0087_[5]),
    .O(s0_data_o[5])
  );
OBUF  _1188_ (
    .I(_0087_[6]),
    .O(s0_data_o[6])
  );
OBUF  _1189_ (
    .I(_0087_[7]),
    .O(s0_data_o[7])
  );
OBUF  _1190_ (
    .I(_0087_[8]),
    .O(s0_data_o[8])
  );
OBUF  _1191_ (
    .I(_0087_[9]),
    .O(s0_data_o[9])
  );
IBUF  _1192_ (
    .I(s0_err_i),
    .O(_0088_)
  );
IBUF  _1193_ (
    .I(s0_rty_i),
    .O(_0089_)
  );
OBUF  _1194_ (
    .I(_0090_[0]),
    .O(s0_sel_o[0])
  );
OBUF  _1195_ (
    .I(_0090_[1]),
    .O(s0_sel_o[1])
  );
OBUF  _1196_ (
    .I(_0090_[2]),
    .O(s0_sel_o[2])
  );
OBUF  _1197_ (
    .I(_0090_[3]),
    .O(s0_sel_o[3])
  );
OBUF  _1198_ (
    .I(_0091_),
    .O(s0_stb_o)
  );
OBUF  _1199_ (
    .I(_0092_),
    .O(s0_we_o)
  );
IBUF  _1200_ (
    .I(s10_ack_i),
    .O(_0093_)
  );
OBUF  _1201_ (
    .I(_0094_[0]),
    .O(s10_addr_o[0])
  );
OBUF  _1202_ (
    .I(_0094_[1]),
    .O(s10_addr_o[1])
  );
OBUF  _1203_ (
    .I(_0094_[10]),
    .O(s10_addr_o[10])
  );
OBUF  _1204_ (
    .I(_0094_[11]),
    .O(s10_addr_o[11])
  );
OBUF  _1205_ (
    .I(_0094_[12]),
    .O(s10_addr_o[12])
  );
OBUF  _1206_ (
    .I(_0094_[13]),
    .O(s10_addr_o[13])
  );
OBUF  _1207_ (
    .I(_0094_[14]),
    .O(s10_addr_o[14])
  );
OBUF  _1208_ (
    .I(_0094_[15]),
    .O(s10_addr_o[15])
  );
OBUF  _1209_ (
    .I(_0094_[16]),
    .O(s10_addr_o[16])
  );
OBUF  _1210_ (
    .I(_0094_[17]),
    .O(s10_addr_o[17])
  );
OBUF  _1211_ (
    .I(_0094_[18]),
    .O(s10_addr_o[18])
  );
OBUF  _1212_ (
    .I(_0094_[19]),
    .O(s10_addr_o[19])
  );
OBUF  _1213_ (
    .I(_0094_[2]),
    .O(s10_addr_o[2])
  );
OBUF  _1214_ (
    .I(_0094_[20]),
    .O(s10_addr_o[20])
  );
OBUF  _1215_ (
    .I(_0094_[21]),
    .O(s10_addr_o[21])
  );
OBUF  _1216_ (
    .I(_0094_[22]),
    .O(s10_addr_o[22])
  );
OBUF  _1217_ (
    .I(_0094_[23]),
    .O(s10_addr_o[23])
  );
OBUF  _1218_ (
    .I(_0094_[24]),
    .O(s10_addr_o[24])
  );
OBUF  _1219_ (
    .I(_0094_[25]),
    .O(s10_addr_o[25])
  );
OBUF  _1220_ (
    .I(_0094_[26]),
    .O(s10_addr_o[26])
  );
OBUF  _1221_ (
    .I(_0094_[27]),
    .O(s10_addr_o[27])
  );
OBUF  _1222_ (
    .I(_0094_[28]),
    .O(s10_addr_o[28])
  );
OBUF  _1223_ (
    .I(_0094_[29]),
    .O(s10_addr_o[29])
  );
OBUF  _1224_ (
    .I(_0094_[3]),
    .O(s10_addr_o[3])
  );
OBUF  _1225_ (
    .I(_0094_[30]),
    .O(s10_addr_o[30])
  );
OBUF  _1226_ (
    .I(_0094_[31]),
    .O(s10_addr_o[31])
  );
OBUF  _1227_ (
    .I(_0094_[4]),
    .O(s10_addr_o[4])
  );
OBUF  _1228_ (
    .I(_0094_[5]),
    .O(s10_addr_o[5])
  );
OBUF  _1229_ (
    .I(_0094_[6]),
    .O(s10_addr_o[6])
  );
OBUF  _1230_ (
    .I(_0094_[7]),
    .O(s10_addr_o[7])
  );
OBUF  _1231_ (
    .I(_0094_[8]),
    .O(s10_addr_o[8])
  );
OBUF  _1232_ (
    .I(_0094_[9]),
    .O(s10_addr_o[9])
  );
OBUF  _1233_ (
    .I(_0095_),
    .O(s10_cyc_o)
  );
IBUF  _1234_ (
    .I(s10_data_i[0]),
    .O(_0096_[0])
  );
IBUF  _1235_ (
    .I(s10_data_i[1]),
    .O(_0096_[1])
  );
IBUF  _1236_ (
    .I(s10_data_i[10]),
    .O(_0096_[10])
  );
IBUF  _1237_ (
    .I(s10_data_i[11]),
    .O(_0096_[11])
  );
IBUF  _1238_ (
    .I(s10_data_i[12]),
    .O(_0096_[12])
  );
IBUF  _1239_ (
    .I(s10_data_i[13]),
    .O(_0096_[13])
  );
IBUF  _1240_ (
    .I(s10_data_i[14]),
    .O(_0096_[14])
  );
IBUF  _1241_ (
    .I(s10_data_i[15]),
    .O(_0096_[15])
  );
IBUF  _1242_ (
    .I(s10_data_i[16]),
    .O(_0096_[16])
  );
IBUF  _1243_ (
    .I(s10_data_i[17]),
    .O(_0096_[17])
  );
IBUF  _1244_ (
    .I(s10_data_i[18]),
    .O(_0096_[18])
  );
IBUF  _1245_ (
    .I(s10_data_i[19]),
    .O(_0096_[19])
  );
IBUF  _1246_ (
    .I(s10_data_i[2]),
    .O(_0096_[2])
  );
IBUF  _1247_ (
    .I(s10_data_i[20]),
    .O(_0096_[20])
  );
IBUF  _1248_ (
    .I(s10_data_i[21]),
    .O(_0096_[21])
  );
IBUF  _1249_ (
    .I(s10_data_i[22]),
    .O(_0096_[22])
  );
IBUF  _1250_ (
    .I(s10_data_i[23]),
    .O(_0096_[23])
  );
IBUF  _1251_ (
    .I(s10_data_i[24]),
    .O(_0096_[24])
  );
IBUF  _1252_ (
    .I(s10_data_i[25]),
    .O(_0096_[25])
  );
IBUF  _1253_ (
    .I(s10_data_i[26]),
    .O(_0096_[26])
  );
IBUF  _1254_ (
    .I(s10_data_i[27]),
    .O(_0096_[27])
  );
IBUF  _1255_ (
    .I(s10_data_i[28]),
    .O(_0096_[28])
  );
IBUF  _1256_ (
    .I(s10_data_i[29]),
    .O(_0096_[29])
  );
IBUF  _1257_ (
    .I(s10_data_i[3]),
    .O(_0096_[3])
  );
IBUF  _1258_ (
    .I(s10_data_i[30]),
    .O(_0096_[30])
  );
IBUF  _1259_ (
    .I(s10_data_i[31]),
    .O(_0096_[31])
  );
IBUF  _1260_ (
    .I(s10_data_i[4]),
    .O(_0096_[4])
  );
IBUF  _1261_ (
    .I(s10_data_i[5]),
    .O(_0096_[5])
  );
IBUF  _1262_ (
    .I(s10_data_i[6]),
    .O(_0096_[6])
  );
IBUF  _1263_ (
    .I(s10_data_i[7]),
    .O(_0096_[7])
  );
IBUF  _1264_ (
    .I(s10_data_i[8]),
    .O(_0096_[8])
  );
IBUF  _1265_ (
    .I(s10_data_i[9]),
    .O(_0096_[9])
  );
OBUF  _1266_ (
    .I(_0097_[0]),
    .O(s10_data_o[0])
  );
OBUF  _1267_ (
    .I(_0097_[1]),
    .O(s10_data_o[1])
  );
OBUF  _1268_ (
    .I(_0097_[10]),
    .O(s10_data_o[10])
  );
OBUF  _1269_ (
    .I(_0097_[11]),
    .O(s10_data_o[11])
  );
OBUF  _1270_ (
    .I(_0097_[12]),
    .O(s10_data_o[12])
  );
OBUF  _1271_ (
    .I(_0097_[13]),
    .O(s10_data_o[13])
  );
OBUF  _1272_ (
    .I(_0097_[14]),
    .O(s10_data_o[14])
  );
OBUF  _1273_ (
    .I(_0097_[15]),
    .O(s10_data_o[15])
  );
OBUF  _1274_ (
    .I(_0097_[16]),
    .O(s10_data_o[16])
  );
OBUF  _1275_ (
    .I(_0097_[17]),
    .O(s10_data_o[17])
  );
OBUF  _1276_ (
    .I(_0097_[18]),
    .O(s10_data_o[18])
  );
OBUF  _1277_ (
    .I(_0097_[19]),
    .O(s10_data_o[19])
  );
OBUF  _1278_ (
    .I(_0097_[2]),
    .O(s10_data_o[2])
  );
OBUF  _1279_ (
    .I(_0097_[20]),
    .O(s10_data_o[20])
  );
OBUF  _1280_ (
    .I(_0097_[21]),
    .O(s10_data_o[21])
  );
OBUF  _1281_ (
    .I(_0097_[22]),
    .O(s10_data_o[22])
  );
OBUF  _1282_ (
    .I(_0097_[23]),
    .O(s10_data_o[23])
  );
OBUF  _1283_ (
    .I(_0097_[24]),
    .O(s10_data_o[24])
  );
OBUF  _1284_ (
    .I(_0097_[25]),
    .O(s10_data_o[25])
  );
OBUF  _1285_ (
    .I(_0097_[26]),
    .O(s10_data_o[26])
  );
OBUF  _1286_ (
    .I(_0097_[27]),
    .O(s10_data_o[27])
  );
OBUF  _1287_ (
    .I(_0097_[28]),
    .O(s10_data_o[28])
  );
OBUF  _1288_ (
    .I(_0097_[29]),
    .O(s10_data_o[29])
  );
OBUF  _1289_ (
    .I(_0097_[3]),
    .O(s10_data_o[3])
  );
OBUF  _1290_ (
    .I(_0097_[30]),
    .O(s10_data_o[30])
  );
OBUF  _1291_ (
    .I(_0097_[31]),
    .O(s10_data_o[31])
  );
OBUF  _1292_ (
    .I(_0097_[4]),
    .O(s10_data_o[4])
  );
OBUF  _1293_ (
    .I(_0097_[5]),
    .O(s10_data_o[5])
  );
OBUF  _1294_ (
    .I(_0097_[6]),
    .O(s10_data_o[6])
  );
OBUF  _1295_ (
    .I(_0097_[7]),
    .O(s10_data_o[7])
  );
OBUF  _1296_ (
    .I(_0097_[8]),
    .O(s10_data_o[8])
  );
OBUF  _1297_ (
    .I(_0097_[9]),
    .O(s10_data_o[9])
  );
IBUF  _1298_ (
    .I(s10_err_i),
    .O(_0098_)
  );
IBUF  _1299_ (
    .I(s10_rty_i),
    .O(_0099_)
  );
OBUF  _1300_ (
    .I(_0100_[0]),
    .O(s10_sel_o[0])
  );
OBUF  _1301_ (
    .I(_0100_[1]),
    .O(s10_sel_o[1])
  );
OBUF  _1302_ (
    .I(_0100_[2]),
    .O(s10_sel_o[2])
  );
OBUF  _1303_ (
    .I(_0100_[3]),
    .O(s10_sel_o[3])
  );
OBUF  _1304_ (
    .I(_0101_),
    .O(s10_stb_o)
  );
OBUF  _1305_ (
    .I(_0102_),
    .O(s10_we_o)
  );
IBUF  _1306_ (
    .I(s11_ack_i),
    .O(_0103_)
  );
OBUF  _1307_ (
    .I(_0104_[0]),
    .O(s11_addr_o[0])
  );
OBUF  _1308_ (
    .I(_0104_[1]),
    .O(s11_addr_o[1])
  );
OBUF  _1309_ (
    .I(_0104_[10]),
    .O(s11_addr_o[10])
  );
OBUF  _1310_ (
    .I(_0104_[11]),
    .O(s11_addr_o[11])
  );
OBUF  _1311_ (
    .I(_0104_[12]),
    .O(s11_addr_o[12])
  );
OBUF  _1312_ (
    .I(_0104_[13]),
    .O(s11_addr_o[13])
  );
OBUF  _1313_ (
    .I(_0104_[14]),
    .O(s11_addr_o[14])
  );
OBUF  _1314_ (
    .I(_0104_[15]),
    .O(s11_addr_o[15])
  );
OBUF  _1315_ (
    .I(_0104_[16]),
    .O(s11_addr_o[16])
  );
OBUF  _1316_ (
    .I(_0104_[17]),
    .O(s11_addr_o[17])
  );
OBUF  _1317_ (
    .I(_0104_[18]),
    .O(s11_addr_o[18])
  );
OBUF  _1318_ (
    .I(_0104_[19]),
    .O(s11_addr_o[19])
  );
OBUF  _1319_ (
    .I(_0104_[2]),
    .O(s11_addr_o[2])
  );
OBUF  _1320_ (
    .I(_0104_[20]),
    .O(s11_addr_o[20])
  );
OBUF  _1321_ (
    .I(_0104_[21]),
    .O(s11_addr_o[21])
  );
OBUF  _1322_ (
    .I(_0104_[22]),
    .O(s11_addr_o[22])
  );
OBUF  _1323_ (
    .I(_0104_[23]),
    .O(s11_addr_o[23])
  );
OBUF  _1324_ (
    .I(_0104_[24]),
    .O(s11_addr_o[24])
  );
OBUF  _1325_ (
    .I(_0104_[25]),
    .O(s11_addr_o[25])
  );
OBUF  _1326_ (
    .I(_0104_[26]),
    .O(s11_addr_o[26])
  );
OBUF  _1327_ (
    .I(_0104_[27]),
    .O(s11_addr_o[27])
  );
OBUF  _1328_ (
    .I(_0104_[28]),
    .O(s11_addr_o[28])
  );
OBUF  _1329_ (
    .I(_0104_[29]),
    .O(s11_addr_o[29])
  );
OBUF  _1330_ (
    .I(_0104_[3]),
    .O(s11_addr_o[3])
  );
OBUF  _1331_ (
    .I(_0104_[30]),
    .O(s11_addr_o[30])
  );
OBUF  _1332_ (
    .I(_0104_[31]),
    .O(s11_addr_o[31])
  );
OBUF  _1333_ (
    .I(_0104_[4]),
    .O(s11_addr_o[4])
  );
OBUF  _1334_ (
    .I(_0104_[5]),
    .O(s11_addr_o[5])
  );
OBUF  _1335_ (
    .I(_0104_[6]),
    .O(s11_addr_o[6])
  );
OBUF  _1336_ (
    .I(_0104_[7]),
    .O(s11_addr_o[7])
  );
OBUF  _1337_ (
    .I(_0104_[8]),
    .O(s11_addr_o[8])
  );
OBUF  _1338_ (
    .I(_0104_[9]),
    .O(s11_addr_o[9])
  );
OBUF  _1339_ (
    .I(_0105_),
    .O(s11_cyc_o)
  );
IBUF  _1340_ (
    .I(s11_data_i[0]),
    .O(_0106_[0])
  );
IBUF  _1341_ (
    .I(s11_data_i[1]),
    .O(_0106_[1])
  );
IBUF  _1342_ (
    .I(s11_data_i[10]),
    .O(_0106_[10])
  );
IBUF  _1343_ (
    .I(s11_data_i[11]),
    .O(_0106_[11])
  );
IBUF  _1344_ (
    .I(s11_data_i[12]),
    .O(_0106_[12])
  );
IBUF  _1345_ (
    .I(s11_data_i[13]),
    .O(_0106_[13])
  );
IBUF  _1346_ (
    .I(s11_data_i[14]),
    .O(_0106_[14])
  );
IBUF  _1347_ (
    .I(s11_data_i[15]),
    .O(_0106_[15])
  );
IBUF  _1348_ (
    .I(s11_data_i[16]),
    .O(_0106_[16])
  );
IBUF  _1349_ (
    .I(s11_data_i[17]),
    .O(_0106_[17])
  );
IBUF  _1350_ (
    .I(s11_data_i[18]),
    .O(_0106_[18])
  );
IBUF  _1351_ (
    .I(s11_data_i[19]),
    .O(_0106_[19])
  );
IBUF  _1352_ (
    .I(s11_data_i[2]),
    .O(_0106_[2])
  );
IBUF  _1353_ (
    .I(s11_data_i[20]),
    .O(_0106_[20])
  );
IBUF  _1354_ (
    .I(s11_data_i[21]),
    .O(_0106_[21])
  );
IBUF  _1355_ (
    .I(s11_data_i[22]),
    .O(_0106_[22])
  );
IBUF  _1356_ (
    .I(s11_data_i[23]),
    .O(_0106_[23])
  );
IBUF  _1357_ (
    .I(s11_data_i[24]),
    .O(_0106_[24])
  );
IBUF  _1358_ (
    .I(s11_data_i[25]),
    .O(_0106_[25])
  );
IBUF  _1359_ (
    .I(s11_data_i[26]),
    .O(_0106_[26])
  );
IBUF  _1360_ (
    .I(s11_data_i[27]),
    .O(_0106_[27])
  );
IBUF  _1361_ (
    .I(s11_data_i[28]),
    .O(_0106_[28])
  );
IBUF  _1362_ (
    .I(s11_data_i[29]),
    .O(_0106_[29])
  );
IBUF  _1363_ (
    .I(s11_data_i[3]),
    .O(_0106_[3])
  );
IBUF  _1364_ (
    .I(s11_data_i[30]),
    .O(_0106_[30])
  );
IBUF  _1365_ (
    .I(s11_data_i[31]),
    .O(_0106_[31])
  );
IBUF  _1366_ (
    .I(s11_data_i[4]),
    .O(_0106_[4])
  );
IBUF  _1367_ (
    .I(s11_data_i[5]),
    .O(_0106_[5])
  );
IBUF  _1368_ (
    .I(s11_data_i[6]),
    .O(_0106_[6])
  );
IBUF  _1369_ (
    .I(s11_data_i[7]),
    .O(_0106_[7])
  );
IBUF  _1370_ (
    .I(s11_data_i[8]),
    .O(_0106_[8])
  );
IBUF  _1371_ (
    .I(s11_data_i[9]),
    .O(_0106_[9])
  );
OBUF  _1372_ (
    .I(_0107_[0]),
    .O(s11_data_o[0])
  );
OBUF  _1373_ (
    .I(_0107_[1]),
    .O(s11_data_o[1])
  );
OBUF  _1374_ (
    .I(_0107_[10]),
    .O(s11_data_o[10])
  );
OBUF  _1375_ (
    .I(_0107_[11]),
    .O(s11_data_o[11])
  );
OBUF  _1376_ (
    .I(_0107_[12]),
    .O(s11_data_o[12])
  );
OBUF  _1377_ (
    .I(_0107_[13]),
    .O(s11_data_o[13])
  );
OBUF  _1378_ (
    .I(_0107_[14]),
    .O(s11_data_o[14])
  );
OBUF  _1379_ (
    .I(_0107_[15]),
    .O(s11_data_o[15])
  );
OBUF  _1380_ (
    .I(_0107_[16]),
    .O(s11_data_o[16])
  );
OBUF  _1381_ (
    .I(_0107_[17]),
    .O(s11_data_o[17])
  );
OBUF  _1382_ (
    .I(_0107_[18]),
    .O(s11_data_o[18])
  );
OBUF  _1383_ (
    .I(_0107_[19]),
    .O(s11_data_o[19])
  );
OBUF  _1384_ (
    .I(_0107_[2]),
    .O(s11_data_o[2])
  );
OBUF  _1385_ (
    .I(_0107_[20]),
    .O(s11_data_o[20])
  );
OBUF  _1386_ (
    .I(_0107_[21]),
    .O(s11_data_o[21])
  );
OBUF  _1387_ (
    .I(_0107_[22]),
    .O(s11_data_o[22])
  );
OBUF  _1388_ (
    .I(_0107_[23]),
    .O(s11_data_o[23])
  );
OBUF  _1389_ (
    .I(_0107_[24]),
    .O(s11_data_o[24])
  );
OBUF  _1390_ (
    .I(_0107_[25]),
    .O(s11_data_o[25])
  );
OBUF  _1391_ (
    .I(_0107_[26]),
    .O(s11_data_o[26])
  );
OBUF  _1392_ (
    .I(_0107_[27]),
    .O(s11_data_o[27])
  );
OBUF  _1393_ (
    .I(_0107_[28]),
    .O(s11_data_o[28])
  );
OBUF  _1394_ (
    .I(_0107_[29]),
    .O(s11_data_o[29])
  );
OBUF  _1395_ (
    .I(_0107_[3]),
    .O(s11_data_o[3])
  );
OBUF  _1396_ (
    .I(_0107_[30]),
    .O(s11_data_o[30])
  );
OBUF  _1397_ (
    .I(_0107_[31]),
    .O(s11_data_o[31])
  );
OBUF  _1398_ (
    .I(_0107_[4]),
    .O(s11_data_o[4])
  );
OBUF  _1399_ (
    .I(_0107_[5]),
    .O(s11_data_o[5])
  );
OBUF  _1400_ (
    .I(_0107_[6]),
    .O(s11_data_o[6])
  );
OBUF  _1401_ (
    .I(_0107_[7]),
    .O(s11_data_o[7])
  );
OBUF  _1402_ (
    .I(_0107_[8]),
    .O(s11_data_o[8])
  );
OBUF  _1403_ (
    .I(_0107_[9]),
    .O(s11_data_o[9])
  );
IBUF  _1404_ (
    .I(s11_err_i),
    .O(_0108_)
  );
IBUF  _1405_ (
    .I(s11_rty_i),
    .O(_0109_)
  );
OBUF  _1406_ (
    .I(_0110_[0]),
    .O(s11_sel_o[0])
  );
OBUF  _1407_ (
    .I(_0110_[1]),
    .O(s11_sel_o[1])
  );
OBUF  _1408_ (
    .I(_0110_[2]),
    .O(s11_sel_o[2])
  );
OBUF  _1409_ (
    .I(_0110_[3]),
    .O(s11_sel_o[3])
  );
OBUF  _1410_ (
    .I(_0111_),
    .O(s11_stb_o)
  );
OBUF  _1411_ (
    .I(_0112_),
    .O(s11_we_o)
  );
IBUF  _1412_ (
    .I(s12_ack_i),
    .O(_0113_)
  );
OBUF  _1413_ (
    .I(_0114_[0]),
    .O(s12_addr_o[0])
  );
OBUF  _1414_ (
    .I(_0114_[1]),
    .O(s12_addr_o[1])
  );
OBUF  _1415_ (
    .I(_0114_[10]),
    .O(s12_addr_o[10])
  );
OBUF  _1416_ (
    .I(_0114_[11]),
    .O(s12_addr_o[11])
  );
OBUF  _1417_ (
    .I(_0114_[12]),
    .O(s12_addr_o[12])
  );
OBUF  _1418_ (
    .I(_0114_[13]),
    .O(s12_addr_o[13])
  );
OBUF  _1419_ (
    .I(_0114_[14]),
    .O(s12_addr_o[14])
  );
OBUF  _1420_ (
    .I(_0114_[15]),
    .O(s12_addr_o[15])
  );
OBUF  _1421_ (
    .I(_0114_[16]),
    .O(s12_addr_o[16])
  );
OBUF  _1422_ (
    .I(_0114_[17]),
    .O(s12_addr_o[17])
  );
OBUF  _1423_ (
    .I(_0114_[18]),
    .O(s12_addr_o[18])
  );
OBUF  _1424_ (
    .I(_0114_[19]),
    .O(s12_addr_o[19])
  );
OBUF  _1425_ (
    .I(_0114_[2]),
    .O(s12_addr_o[2])
  );
OBUF  _1426_ (
    .I(_0114_[20]),
    .O(s12_addr_o[20])
  );
OBUF  _1427_ (
    .I(_0114_[21]),
    .O(s12_addr_o[21])
  );
OBUF  _1428_ (
    .I(_0114_[22]),
    .O(s12_addr_o[22])
  );
OBUF  _1429_ (
    .I(_0114_[23]),
    .O(s12_addr_o[23])
  );
OBUF  _1430_ (
    .I(_0114_[24]),
    .O(s12_addr_o[24])
  );
OBUF  _1431_ (
    .I(_0114_[25]),
    .O(s12_addr_o[25])
  );
OBUF  _1432_ (
    .I(_0114_[26]),
    .O(s12_addr_o[26])
  );
OBUF  _1433_ (
    .I(_0114_[27]),
    .O(s12_addr_o[27])
  );
OBUF  _1434_ (
    .I(_0114_[28]),
    .O(s12_addr_o[28])
  );
OBUF  _1435_ (
    .I(_0114_[29]),
    .O(s12_addr_o[29])
  );
OBUF  _1436_ (
    .I(_0114_[3]),
    .O(s12_addr_o[3])
  );
OBUF  _1437_ (
    .I(_0114_[30]),
    .O(s12_addr_o[30])
  );
OBUF  _1438_ (
    .I(_0114_[31]),
    .O(s12_addr_o[31])
  );
OBUF  _1439_ (
    .I(_0114_[4]),
    .O(s12_addr_o[4])
  );
OBUF  _1440_ (
    .I(_0114_[5]),
    .O(s12_addr_o[5])
  );
OBUF  _1441_ (
    .I(_0114_[6]),
    .O(s12_addr_o[6])
  );
OBUF  _1442_ (
    .I(_0114_[7]),
    .O(s12_addr_o[7])
  );
OBUF  _1443_ (
    .I(_0114_[8]),
    .O(s12_addr_o[8])
  );
OBUF  _1444_ (
    .I(_0114_[9]),
    .O(s12_addr_o[9])
  );
OBUF  _1445_ (
    .I(_0115_),
    .O(s12_cyc_o)
  );
IBUF  _1446_ (
    .I(s12_data_i[0]),
    .O(_0116_[0])
  );
IBUF  _1447_ (
    .I(s12_data_i[1]),
    .O(_0116_[1])
  );
IBUF  _1448_ (
    .I(s12_data_i[10]),
    .O(_0116_[10])
  );
IBUF  _1449_ (
    .I(s12_data_i[11]),
    .O(_0116_[11])
  );
IBUF  _1450_ (
    .I(s12_data_i[12]),
    .O(_0116_[12])
  );
IBUF  _1451_ (
    .I(s12_data_i[13]),
    .O(_0116_[13])
  );
IBUF  _1452_ (
    .I(s12_data_i[14]),
    .O(_0116_[14])
  );
IBUF  _1453_ (
    .I(s12_data_i[15]),
    .O(_0116_[15])
  );
IBUF  _1454_ (
    .I(s12_data_i[16]),
    .O(_0116_[16])
  );
IBUF  _1455_ (
    .I(s12_data_i[17]),
    .O(_0116_[17])
  );
IBUF  _1456_ (
    .I(s12_data_i[18]),
    .O(_0116_[18])
  );
IBUF  _1457_ (
    .I(s12_data_i[19]),
    .O(_0116_[19])
  );
IBUF  _1458_ (
    .I(s12_data_i[2]),
    .O(_0116_[2])
  );
IBUF  _1459_ (
    .I(s12_data_i[20]),
    .O(_0116_[20])
  );
IBUF  _1460_ (
    .I(s12_data_i[21]),
    .O(_0116_[21])
  );
IBUF  _1461_ (
    .I(s12_data_i[22]),
    .O(_0116_[22])
  );
IBUF  _1462_ (
    .I(s12_data_i[23]),
    .O(_0116_[23])
  );
IBUF  _1463_ (
    .I(s12_data_i[24]),
    .O(_0116_[24])
  );
IBUF  _1464_ (
    .I(s12_data_i[25]),
    .O(_0116_[25])
  );
IBUF  _1465_ (
    .I(s12_data_i[26]),
    .O(_0116_[26])
  );
IBUF  _1466_ (
    .I(s12_data_i[27]),
    .O(_0116_[27])
  );
IBUF  _1467_ (
    .I(s12_data_i[28]),
    .O(_0116_[28])
  );
IBUF  _1468_ (
    .I(s12_data_i[29]),
    .O(_0116_[29])
  );
IBUF  _1469_ (
    .I(s12_data_i[3]),
    .O(_0116_[3])
  );
IBUF  _1470_ (
    .I(s12_data_i[30]),
    .O(_0116_[30])
  );
IBUF  _1471_ (
    .I(s12_data_i[31]),
    .O(_0116_[31])
  );
IBUF  _1472_ (
    .I(s12_data_i[4]),
    .O(_0116_[4])
  );
IBUF  _1473_ (
    .I(s12_data_i[5]),
    .O(_0116_[5])
  );
IBUF  _1474_ (
    .I(s12_data_i[6]),
    .O(_0116_[6])
  );
IBUF  _1475_ (
    .I(s12_data_i[7]),
    .O(_0116_[7])
  );
IBUF  _1476_ (
    .I(s12_data_i[8]),
    .O(_0116_[8])
  );
IBUF  _1477_ (
    .I(s12_data_i[9]),
    .O(_0116_[9])
  );
OBUF  _1478_ (
    .I(_0117_[0]),
    .O(s12_data_o[0])
  );
OBUF  _1479_ (
    .I(_0117_[1]),
    .O(s12_data_o[1])
  );
OBUF  _1480_ (
    .I(_0117_[10]),
    .O(s12_data_o[10])
  );
OBUF  _1481_ (
    .I(_0117_[11]),
    .O(s12_data_o[11])
  );
OBUF  _1482_ (
    .I(_0117_[12]),
    .O(s12_data_o[12])
  );
OBUF  _1483_ (
    .I(_0117_[13]),
    .O(s12_data_o[13])
  );
OBUF  _1484_ (
    .I(_0117_[14]),
    .O(s12_data_o[14])
  );
OBUF  _1485_ (
    .I(_0117_[15]),
    .O(s12_data_o[15])
  );
OBUF  _1486_ (
    .I(_0117_[16]),
    .O(s12_data_o[16])
  );
OBUF  _1487_ (
    .I(_0117_[17]),
    .O(s12_data_o[17])
  );
OBUF  _1488_ (
    .I(_0117_[18]),
    .O(s12_data_o[18])
  );
OBUF  _1489_ (
    .I(_0117_[19]),
    .O(s12_data_o[19])
  );
OBUF  _1490_ (
    .I(_0117_[2]),
    .O(s12_data_o[2])
  );
OBUF  _1491_ (
    .I(_0117_[20]),
    .O(s12_data_o[20])
  );
OBUF  _1492_ (
    .I(_0117_[21]),
    .O(s12_data_o[21])
  );
OBUF  _1493_ (
    .I(_0117_[22]),
    .O(s12_data_o[22])
  );
OBUF  _1494_ (
    .I(_0117_[23]),
    .O(s12_data_o[23])
  );
OBUF  _1495_ (
    .I(_0117_[24]),
    .O(s12_data_o[24])
  );
OBUF  _1496_ (
    .I(_0117_[25]),
    .O(s12_data_o[25])
  );
OBUF  _1497_ (
    .I(_0117_[26]),
    .O(s12_data_o[26])
  );
OBUF  _1498_ (
    .I(_0117_[27]),
    .O(s12_data_o[27])
  );
OBUF  _1499_ (
    .I(_0117_[28]),
    .O(s12_data_o[28])
  );
OBUF  _1500_ (
    .I(_0117_[29]),
    .O(s12_data_o[29])
  );
OBUF  _1501_ (
    .I(_0117_[3]),
    .O(s12_data_o[3])
  );
OBUF  _1502_ (
    .I(_0117_[30]),
    .O(s12_data_o[30])
  );
OBUF  _1503_ (
    .I(_0117_[31]),
    .O(s12_data_o[31])
  );
OBUF  _1504_ (
    .I(_0117_[4]),
    .O(s12_data_o[4])
  );
OBUF  _1505_ (
    .I(_0117_[5]),
    .O(s12_data_o[5])
  );
OBUF  _1506_ (
    .I(_0117_[6]),
    .O(s12_data_o[6])
  );
OBUF  _1507_ (
    .I(_0117_[7]),
    .O(s12_data_o[7])
  );
OBUF  _1508_ (
    .I(_0117_[8]),
    .O(s12_data_o[8])
  );
OBUF  _1509_ (
    .I(_0117_[9]),
    .O(s12_data_o[9])
  );
IBUF  _1510_ (
    .I(s12_err_i),
    .O(_0118_)
  );
IBUF  _1511_ (
    .I(s12_rty_i),
    .O(_0119_)
  );
OBUF  _1512_ (
    .I(_0120_[0]),
    .O(s12_sel_o[0])
  );
OBUF  _1513_ (
    .I(_0120_[1]),
    .O(s12_sel_o[1])
  );
OBUF  _1514_ (
    .I(_0120_[2]),
    .O(s12_sel_o[2])
  );
OBUF  _1515_ (
    .I(_0120_[3]),
    .O(s12_sel_o[3])
  );
OBUF  _1516_ (
    .I(_0121_),
    .O(s12_stb_o)
  );
OBUF  _1517_ (
    .I(_0122_),
    .O(s12_we_o)
  );
IBUF  _1518_ (
    .I(s13_ack_i),
    .O(_0123_)
  );
OBUF  _1519_ (
    .I(_0124_[0]),
    .O(s13_addr_o[0])
  );
OBUF  _1520_ (
    .I(_0124_[1]),
    .O(s13_addr_o[1])
  );
OBUF  _1521_ (
    .I(_0124_[10]),
    .O(s13_addr_o[10])
  );
OBUF  _1522_ (
    .I(_0124_[11]),
    .O(s13_addr_o[11])
  );
OBUF  _1523_ (
    .I(_0124_[12]),
    .O(s13_addr_o[12])
  );
OBUF  _1524_ (
    .I(_0124_[13]),
    .O(s13_addr_o[13])
  );
OBUF  _1525_ (
    .I(_0124_[14]),
    .O(s13_addr_o[14])
  );
OBUF  _1526_ (
    .I(_0124_[15]),
    .O(s13_addr_o[15])
  );
OBUF  _1527_ (
    .I(_0124_[16]),
    .O(s13_addr_o[16])
  );
OBUF  _1528_ (
    .I(_0124_[17]),
    .O(s13_addr_o[17])
  );
OBUF  _1529_ (
    .I(_0124_[18]),
    .O(s13_addr_o[18])
  );
OBUF  _1530_ (
    .I(_0124_[19]),
    .O(s13_addr_o[19])
  );
OBUF  _1531_ (
    .I(_0124_[2]),
    .O(s13_addr_o[2])
  );
OBUF  _1532_ (
    .I(_0124_[20]),
    .O(s13_addr_o[20])
  );
OBUF  _1533_ (
    .I(_0124_[21]),
    .O(s13_addr_o[21])
  );
OBUF  _1534_ (
    .I(_0124_[22]),
    .O(s13_addr_o[22])
  );
OBUF  _1535_ (
    .I(_0124_[23]),
    .O(s13_addr_o[23])
  );
OBUF  _1536_ (
    .I(_0124_[24]),
    .O(s13_addr_o[24])
  );
OBUF  _1537_ (
    .I(_0124_[25]),
    .O(s13_addr_o[25])
  );
OBUF  _1538_ (
    .I(_0124_[26]),
    .O(s13_addr_o[26])
  );
OBUF  _1539_ (
    .I(_0124_[27]),
    .O(s13_addr_o[27])
  );
OBUF  _1540_ (
    .I(_0124_[28]),
    .O(s13_addr_o[28])
  );
OBUF  _1541_ (
    .I(_0124_[29]),
    .O(s13_addr_o[29])
  );
OBUF  _1542_ (
    .I(_0124_[3]),
    .O(s13_addr_o[3])
  );
OBUF  _1543_ (
    .I(_0124_[30]),
    .O(s13_addr_o[30])
  );
OBUF  _1544_ (
    .I(_0124_[31]),
    .O(s13_addr_o[31])
  );
OBUF  _1545_ (
    .I(_0124_[4]),
    .O(s13_addr_o[4])
  );
OBUF  _1546_ (
    .I(_0124_[5]),
    .O(s13_addr_o[5])
  );
OBUF  _1547_ (
    .I(_0124_[6]),
    .O(s13_addr_o[6])
  );
OBUF  _1548_ (
    .I(_0124_[7]),
    .O(s13_addr_o[7])
  );
OBUF  _1549_ (
    .I(_0124_[8]),
    .O(s13_addr_o[8])
  );
OBUF  _1550_ (
    .I(_0124_[9]),
    .O(s13_addr_o[9])
  );
OBUF  _1551_ (
    .I(_0125_),
    .O(s13_cyc_o)
  );
IBUF  _1552_ (
    .I(s13_data_i[0]),
    .O(_0126_[0])
  );
IBUF  _1553_ (
    .I(s13_data_i[1]),
    .O(_0126_[1])
  );
IBUF  _1554_ (
    .I(s13_data_i[10]),
    .O(_0126_[10])
  );
IBUF  _1555_ (
    .I(s13_data_i[11]),
    .O(_0126_[11])
  );
IBUF  _1556_ (
    .I(s13_data_i[12]),
    .O(_0126_[12])
  );
IBUF  _1557_ (
    .I(s13_data_i[13]),
    .O(_0126_[13])
  );
IBUF  _1558_ (
    .I(s13_data_i[14]),
    .O(_0126_[14])
  );
IBUF  _1559_ (
    .I(s13_data_i[15]),
    .O(_0126_[15])
  );
IBUF  _1560_ (
    .I(s13_data_i[16]),
    .O(_0126_[16])
  );
IBUF  _1561_ (
    .I(s13_data_i[17]),
    .O(_0126_[17])
  );
IBUF  _1562_ (
    .I(s13_data_i[18]),
    .O(_0126_[18])
  );
IBUF  _1563_ (
    .I(s13_data_i[19]),
    .O(_0126_[19])
  );
IBUF  _1564_ (
    .I(s13_data_i[2]),
    .O(_0126_[2])
  );
IBUF  _1565_ (
    .I(s13_data_i[20]),
    .O(_0126_[20])
  );
IBUF  _1566_ (
    .I(s13_data_i[21]),
    .O(_0126_[21])
  );
IBUF  _1567_ (
    .I(s13_data_i[22]),
    .O(_0126_[22])
  );
IBUF  _1568_ (
    .I(s13_data_i[23]),
    .O(_0126_[23])
  );
IBUF  _1569_ (
    .I(s13_data_i[24]),
    .O(_0126_[24])
  );
IBUF  _1570_ (
    .I(s13_data_i[25]),
    .O(_0126_[25])
  );
IBUF  _1571_ (
    .I(s13_data_i[26]),
    .O(_0126_[26])
  );
IBUF  _1572_ (
    .I(s13_data_i[27]),
    .O(_0126_[27])
  );
IBUF  _1573_ (
    .I(s13_data_i[28]),
    .O(_0126_[28])
  );
IBUF  _1574_ (
    .I(s13_data_i[29]),
    .O(_0126_[29])
  );
IBUF  _1575_ (
    .I(s13_data_i[3]),
    .O(_0126_[3])
  );
IBUF  _1576_ (
    .I(s13_data_i[30]),
    .O(_0126_[30])
  );
IBUF  _1577_ (
    .I(s13_data_i[31]),
    .O(_0126_[31])
  );
IBUF  _1578_ (
    .I(s13_data_i[4]),
    .O(_0126_[4])
  );
IBUF  _1579_ (
    .I(s13_data_i[5]),
    .O(_0126_[5])
  );
IBUF  _1580_ (
    .I(s13_data_i[6]),
    .O(_0126_[6])
  );
IBUF  _1581_ (
    .I(s13_data_i[7]),
    .O(_0126_[7])
  );
IBUF  _1582_ (
    .I(s13_data_i[8]),
    .O(_0126_[8])
  );
IBUF  _1583_ (
    .I(s13_data_i[9]),
    .O(_0126_[9])
  );
OBUF  _1584_ (
    .I(_0127_[0]),
    .O(s13_data_o[0])
  );
OBUF  _1585_ (
    .I(_0127_[1]),
    .O(s13_data_o[1])
  );
OBUF  _1586_ (
    .I(_0127_[10]),
    .O(s13_data_o[10])
  );
OBUF  _1587_ (
    .I(_0127_[11]),
    .O(s13_data_o[11])
  );
OBUF  _1588_ (
    .I(_0127_[12]),
    .O(s13_data_o[12])
  );
OBUF  _1589_ (
    .I(_0127_[13]),
    .O(s13_data_o[13])
  );
OBUF  _1590_ (
    .I(_0127_[14]),
    .O(s13_data_o[14])
  );
OBUF  _1591_ (
    .I(_0127_[15]),
    .O(s13_data_o[15])
  );
OBUF  _1592_ (
    .I(_0127_[16]),
    .O(s13_data_o[16])
  );
OBUF  _1593_ (
    .I(_0127_[17]),
    .O(s13_data_o[17])
  );
OBUF  _1594_ (
    .I(_0127_[18]),
    .O(s13_data_o[18])
  );
OBUF  _1595_ (
    .I(_0127_[19]),
    .O(s13_data_o[19])
  );
OBUF  _1596_ (
    .I(_0127_[2]),
    .O(s13_data_o[2])
  );
OBUF  _1597_ (
    .I(_0127_[20]),
    .O(s13_data_o[20])
  );
OBUF  _1598_ (
    .I(_0127_[21]),
    .O(s13_data_o[21])
  );
OBUF  _1599_ (
    .I(_0127_[22]),
    .O(s13_data_o[22])
  );
OBUF  _1600_ (
    .I(_0127_[23]),
    .O(s13_data_o[23])
  );
OBUF  _1601_ (
    .I(_0127_[24]),
    .O(s13_data_o[24])
  );
OBUF  _1602_ (
    .I(_0127_[25]),
    .O(s13_data_o[25])
  );
OBUF  _1603_ (
    .I(_0127_[26]),
    .O(s13_data_o[26])
  );
OBUF  _1604_ (
    .I(_0127_[27]),
    .O(s13_data_o[27])
  );
OBUF  _1605_ (
    .I(_0127_[28]),
    .O(s13_data_o[28])
  );
OBUF  _1606_ (
    .I(_0127_[29]),
    .O(s13_data_o[29])
  );
OBUF  _1607_ (
    .I(_0127_[3]),
    .O(s13_data_o[3])
  );
OBUF  _1608_ (
    .I(_0127_[30]),
    .O(s13_data_o[30])
  );
OBUF  _1609_ (
    .I(_0127_[31]),
    .O(s13_data_o[31])
  );
OBUF  _1610_ (
    .I(_0127_[4]),
    .O(s13_data_o[4])
  );
OBUF  _1611_ (
    .I(_0127_[5]),
    .O(s13_data_o[5])
  );
OBUF  _1612_ (
    .I(_0127_[6]),
    .O(s13_data_o[6])
  );
OBUF  _1613_ (
    .I(_0127_[7]),
    .O(s13_data_o[7])
  );
OBUF  _1614_ (
    .I(_0127_[8]),
    .O(s13_data_o[8])
  );
OBUF  _1615_ (
    .I(_0127_[9]),
    .O(s13_data_o[9])
  );
IBUF  _1616_ (
    .I(s13_err_i),
    .O(_0128_)
  );
IBUF  _1617_ (
    .I(s13_rty_i),
    .O(_0129_)
  );
OBUF  _1618_ (
    .I(_0130_[0]),
    .O(s13_sel_o[0])
  );
OBUF  _1619_ (
    .I(_0130_[1]),
    .O(s13_sel_o[1])
  );
OBUF  _1620_ (
    .I(_0130_[2]),
    .O(s13_sel_o[2])
  );
OBUF  _1621_ (
    .I(_0130_[3]),
    .O(s13_sel_o[3])
  );
OBUF  _1622_ (
    .I(_0131_),
    .O(s13_stb_o)
  );
OBUF  _1623_ (
    .I(_0132_),
    .O(s13_we_o)
  );
IBUF  _1624_ (
    .I(s14_ack_i),
    .O(_0133_)
  );
OBUF  _1625_ (
    .I(_0134_[0]),
    .O(s14_addr_o[0])
  );
OBUF  _1626_ (
    .I(_0134_[1]),
    .O(s14_addr_o[1])
  );
OBUF  _1627_ (
    .I(_0134_[10]),
    .O(s14_addr_o[10])
  );
OBUF  _1628_ (
    .I(_0134_[11]),
    .O(s14_addr_o[11])
  );
OBUF  _1629_ (
    .I(_0134_[12]),
    .O(s14_addr_o[12])
  );
OBUF  _1630_ (
    .I(_0134_[13]),
    .O(s14_addr_o[13])
  );
OBUF  _1631_ (
    .I(_0134_[14]),
    .O(s14_addr_o[14])
  );
OBUF  _1632_ (
    .I(_0134_[15]),
    .O(s14_addr_o[15])
  );
OBUF  _1633_ (
    .I(_0134_[16]),
    .O(s14_addr_o[16])
  );
OBUF  _1634_ (
    .I(_0134_[17]),
    .O(s14_addr_o[17])
  );
OBUF  _1635_ (
    .I(_0134_[18]),
    .O(s14_addr_o[18])
  );
OBUF  _1636_ (
    .I(_0134_[19]),
    .O(s14_addr_o[19])
  );
OBUF  _1637_ (
    .I(_0134_[2]),
    .O(s14_addr_o[2])
  );
OBUF  _1638_ (
    .I(_0134_[20]),
    .O(s14_addr_o[20])
  );
OBUF  _1639_ (
    .I(_0134_[21]),
    .O(s14_addr_o[21])
  );
OBUF  _1640_ (
    .I(_0134_[22]),
    .O(s14_addr_o[22])
  );
OBUF  _1641_ (
    .I(_0134_[23]),
    .O(s14_addr_o[23])
  );
OBUF  _1642_ (
    .I(_0134_[24]),
    .O(s14_addr_o[24])
  );
OBUF  _1643_ (
    .I(_0134_[25]),
    .O(s14_addr_o[25])
  );
OBUF  _1644_ (
    .I(_0134_[26]),
    .O(s14_addr_o[26])
  );
OBUF  _1645_ (
    .I(_0134_[27]),
    .O(s14_addr_o[27])
  );
OBUF  _1646_ (
    .I(_0134_[28]),
    .O(s14_addr_o[28])
  );
OBUF  _1647_ (
    .I(_0134_[29]),
    .O(s14_addr_o[29])
  );
OBUF  _1648_ (
    .I(_0134_[3]),
    .O(s14_addr_o[3])
  );
OBUF  _1649_ (
    .I(_0134_[30]),
    .O(s14_addr_o[30])
  );
OBUF  _1650_ (
    .I(_0134_[31]),
    .O(s14_addr_o[31])
  );
OBUF  _1651_ (
    .I(_0134_[4]),
    .O(s14_addr_o[4])
  );
OBUF  _1652_ (
    .I(_0134_[5]),
    .O(s14_addr_o[5])
  );
OBUF  _1653_ (
    .I(_0134_[6]),
    .O(s14_addr_o[6])
  );
OBUF  _1654_ (
    .I(_0134_[7]),
    .O(s14_addr_o[7])
  );
OBUF  _1655_ (
    .I(_0134_[8]),
    .O(s14_addr_o[8])
  );
OBUF  _1656_ (
    .I(_0134_[9]),
    .O(s14_addr_o[9])
  );
OBUF  _1657_ (
    .I(_0135_),
    .O(s14_cyc_o)
  );
IBUF  _1658_ (
    .I(s14_data_i[0]),
    .O(_0136_[0])
  );
IBUF  _1659_ (
    .I(s14_data_i[1]),
    .O(_0136_[1])
  );
IBUF  _1660_ (
    .I(s14_data_i[10]),
    .O(_0136_[10])
  );
IBUF  _1661_ (
    .I(s14_data_i[11]),
    .O(_0136_[11])
  );
IBUF  _1662_ (
    .I(s14_data_i[12]),
    .O(_0136_[12])
  );
IBUF  _1663_ (
    .I(s14_data_i[13]),
    .O(_0136_[13])
  );
IBUF  _1664_ (
    .I(s14_data_i[14]),
    .O(_0136_[14])
  );
IBUF  _1665_ (
    .I(s14_data_i[15]),
    .O(_0136_[15])
  );
IBUF  _1666_ (
    .I(s14_data_i[16]),
    .O(_0136_[16])
  );
IBUF  _1667_ (
    .I(s14_data_i[17]),
    .O(_0136_[17])
  );
IBUF  _1668_ (
    .I(s14_data_i[18]),
    .O(_0136_[18])
  );
IBUF  _1669_ (
    .I(s14_data_i[19]),
    .O(_0136_[19])
  );
IBUF  _1670_ (
    .I(s14_data_i[2]),
    .O(_0136_[2])
  );
IBUF  _1671_ (
    .I(s14_data_i[20]),
    .O(_0136_[20])
  );
IBUF  _1672_ (
    .I(s14_data_i[21]),
    .O(_0136_[21])
  );
IBUF  _1673_ (
    .I(s14_data_i[22]),
    .O(_0136_[22])
  );
IBUF  _1674_ (
    .I(s14_data_i[23]),
    .O(_0136_[23])
  );
IBUF  _1675_ (
    .I(s14_data_i[24]),
    .O(_0136_[24])
  );
IBUF  _1676_ (
    .I(s14_data_i[25]),
    .O(_0136_[25])
  );
IBUF  _1677_ (
    .I(s14_data_i[26]),
    .O(_0136_[26])
  );
IBUF  _1678_ (
    .I(s14_data_i[27]),
    .O(_0136_[27])
  );
IBUF  _1679_ (
    .I(s14_data_i[28]),
    .O(_0136_[28])
  );
IBUF  _1680_ (
    .I(s14_data_i[29]),
    .O(_0136_[29])
  );
IBUF  _1681_ (
    .I(s14_data_i[3]),
    .O(_0136_[3])
  );
IBUF  _1682_ (
    .I(s14_data_i[30]),
    .O(_0136_[30])
  );
IBUF  _1683_ (
    .I(s14_data_i[31]),
    .O(_0136_[31])
  );
IBUF  _1684_ (
    .I(s14_data_i[4]),
    .O(_0136_[4])
  );
IBUF  _1685_ (
    .I(s14_data_i[5]),
    .O(_0136_[5])
  );
IBUF  _1686_ (
    .I(s14_data_i[6]),
    .O(_0136_[6])
  );
IBUF  _1687_ (
    .I(s14_data_i[7]),
    .O(_0136_[7])
  );
IBUF  _1688_ (
    .I(s14_data_i[8]),
    .O(_0136_[8])
  );
IBUF  _1689_ (
    .I(s14_data_i[9]),
    .O(_0136_[9])
  );
OBUF  _1690_ (
    .I(_0137_[0]),
    .O(s14_data_o[0])
  );
OBUF  _1691_ (
    .I(_0137_[1]),
    .O(s14_data_o[1])
  );
OBUF  _1692_ (
    .I(_0137_[10]),
    .O(s14_data_o[10])
  );
OBUF  _1693_ (
    .I(_0137_[11]),
    .O(s14_data_o[11])
  );
OBUF  _1694_ (
    .I(_0137_[12]),
    .O(s14_data_o[12])
  );
OBUF  _1695_ (
    .I(_0137_[13]),
    .O(s14_data_o[13])
  );
OBUF  _1696_ (
    .I(_0137_[14]),
    .O(s14_data_o[14])
  );
OBUF  _1697_ (
    .I(_0137_[15]),
    .O(s14_data_o[15])
  );
OBUF  _1698_ (
    .I(_0137_[16]),
    .O(s14_data_o[16])
  );
OBUF  _1699_ (
    .I(_0137_[17]),
    .O(s14_data_o[17])
  );
OBUF  _1700_ (
    .I(_0137_[18]),
    .O(s14_data_o[18])
  );
OBUF  _1701_ (
    .I(_0137_[19]),
    .O(s14_data_o[19])
  );
OBUF  _1702_ (
    .I(_0137_[2]),
    .O(s14_data_o[2])
  );
OBUF  _1703_ (
    .I(_0137_[20]),
    .O(s14_data_o[20])
  );
OBUF  _1704_ (
    .I(_0137_[21]),
    .O(s14_data_o[21])
  );
OBUF  _1705_ (
    .I(_0137_[22]),
    .O(s14_data_o[22])
  );
OBUF  _1706_ (
    .I(_0137_[23]),
    .O(s14_data_o[23])
  );
OBUF  _1707_ (
    .I(_0137_[24]),
    .O(s14_data_o[24])
  );
OBUF  _1708_ (
    .I(_0137_[25]),
    .O(s14_data_o[25])
  );
OBUF  _1709_ (
    .I(_0137_[26]),
    .O(s14_data_o[26])
  );
OBUF  _1710_ (
    .I(_0137_[27]),
    .O(s14_data_o[27])
  );
OBUF  _1711_ (
    .I(_0137_[28]),
    .O(s14_data_o[28])
  );
OBUF  _1712_ (
    .I(_0137_[29]),
    .O(s14_data_o[29])
  );
OBUF  _1713_ (
    .I(_0137_[3]),
    .O(s14_data_o[3])
  );
OBUF  _1714_ (
    .I(_0137_[30]),
    .O(s14_data_o[30])
  );
OBUF  _1715_ (
    .I(_0137_[31]),
    .O(s14_data_o[31])
  );
OBUF  _1716_ (
    .I(_0137_[4]),
    .O(s14_data_o[4])
  );
OBUF  _1717_ (
    .I(_0137_[5]),
    .O(s14_data_o[5])
  );
OBUF  _1718_ (
    .I(_0137_[6]),
    .O(s14_data_o[6])
  );
OBUF  _1719_ (
    .I(_0137_[7]),
    .O(s14_data_o[7])
  );
OBUF  _1720_ (
    .I(_0137_[8]),
    .O(s14_data_o[8])
  );
OBUF  _1721_ (
    .I(_0137_[9]),
    .O(s14_data_o[9])
  );
IBUF  _1722_ (
    .I(s14_err_i),
    .O(_0138_)
  );
IBUF  _1723_ (
    .I(s14_rty_i),
    .O(_0139_)
  );
OBUF  _1724_ (
    .I(_0140_[0]),
    .O(s14_sel_o[0])
  );
OBUF  _1725_ (
    .I(_0140_[1]),
    .O(s14_sel_o[1])
  );
OBUF  _1726_ (
    .I(_0140_[2]),
    .O(s14_sel_o[2])
  );
OBUF  _1727_ (
    .I(_0140_[3]),
    .O(s14_sel_o[3])
  );
OBUF  _1728_ (
    .I(_0141_),
    .O(s14_stb_o)
  );
OBUF  _1729_ (
    .I(_0142_),
    .O(s14_we_o)
  );
IBUF  _1730_ (
    .I(s15_ack_i),
    .O(_0143_)
  );
OBUF  _1731_ (
    .I(_0144_[0]),
    .O(s15_addr_o[0])
  );
OBUF  _1732_ (
    .I(_0144_[1]),
    .O(s15_addr_o[1])
  );
OBUF  _1733_ (
    .I(_0144_[10]),
    .O(s15_addr_o[10])
  );
OBUF  _1734_ (
    .I(_0144_[11]),
    .O(s15_addr_o[11])
  );
OBUF  _1735_ (
    .I(_0144_[12]),
    .O(s15_addr_o[12])
  );
OBUF  _1736_ (
    .I(_0144_[13]),
    .O(s15_addr_o[13])
  );
OBUF  _1737_ (
    .I(_0144_[14]),
    .O(s15_addr_o[14])
  );
OBUF  _1738_ (
    .I(_0144_[15]),
    .O(s15_addr_o[15])
  );
OBUF  _1739_ (
    .I(_0144_[16]),
    .O(s15_addr_o[16])
  );
OBUF  _1740_ (
    .I(_0144_[17]),
    .O(s15_addr_o[17])
  );
OBUF  _1741_ (
    .I(_0144_[18]),
    .O(s15_addr_o[18])
  );
OBUF  _1742_ (
    .I(_0144_[19]),
    .O(s15_addr_o[19])
  );
OBUF  _1743_ (
    .I(_0144_[2]),
    .O(s15_addr_o[2])
  );
OBUF  _1744_ (
    .I(_0144_[20]),
    .O(s15_addr_o[20])
  );
OBUF  _1745_ (
    .I(_0144_[21]),
    .O(s15_addr_o[21])
  );
OBUF  _1746_ (
    .I(_0144_[22]),
    .O(s15_addr_o[22])
  );
OBUF  _1747_ (
    .I(_0144_[23]),
    .O(s15_addr_o[23])
  );
OBUF  _1748_ (
    .I(_0144_[24]),
    .O(s15_addr_o[24])
  );
OBUF  _1749_ (
    .I(_0144_[25]),
    .O(s15_addr_o[25])
  );
OBUF  _1750_ (
    .I(_0144_[26]),
    .O(s15_addr_o[26])
  );
OBUF  _1751_ (
    .I(_0144_[27]),
    .O(s15_addr_o[27])
  );
OBUF  _1752_ (
    .I(_0144_[28]),
    .O(s15_addr_o[28])
  );
OBUF  _1753_ (
    .I(_0144_[29]),
    .O(s15_addr_o[29])
  );
OBUF  _1754_ (
    .I(_0144_[3]),
    .O(s15_addr_o[3])
  );
OBUF  _1755_ (
    .I(_0144_[30]),
    .O(s15_addr_o[30])
  );
OBUF  _1756_ (
    .I(_0144_[31]),
    .O(s15_addr_o[31])
  );
OBUF  _1757_ (
    .I(_0144_[4]),
    .O(s15_addr_o[4])
  );
OBUF  _1758_ (
    .I(_0144_[5]),
    .O(s15_addr_o[5])
  );
OBUF  _1759_ (
    .I(_0144_[6]),
    .O(s15_addr_o[6])
  );
OBUF  _1760_ (
    .I(_0144_[7]),
    .O(s15_addr_o[7])
  );
OBUF  _1761_ (
    .I(_0144_[8]),
    .O(s15_addr_o[8])
  );
OBUF  _1762_ (
    .I(_0144_[9]),
    .O(s15_addr_o[9])
  );
OBUF  _1763_ (
    .I(_0145_),
    .O(s15_cyc_o)
  );
IBUF  _1764_ (
    .I(s15_data_i[0]),
    .O(_0146_[0])
  );
IBUF  _1765_ (
    .I(s15_data_i[1]),
    .O(_0146_[1])
  );
IBUF  _1766_ (
    .I(s15_data_i[10]),
    .O(_0146_[10])
  );
IBUF  _1767_ (
    .I(s15_data_i[11]),
    .O(_0146_[11])
  );
IBUF  _1768_ (
    .I(s15_data_i[12]),
    .O(_0146_[12])
  );
IBUF  _1769_ (
    .I(s15_data_i[13]),
    .O(_0146_[13])
  );
IBUF  _1770_ (
    .I(s15_data_i[14]),
    .O(_0146_[14])
  );
IBUF  _1771_ (
    .I(s15_data_i[15]),
    .O(_0146_[15])
  );
IBUF  _1772_ (
    .I(s15_data_i[16]),
    .O(_0146_[16])
  );
IBUF  _1773_ (
    .I(s15_data_i[17]),
    .O(_0146_[17])
  );
IBUF  _1774_ (
    .I(s15_data_i[18]),
    .O(_0146_[18])
  );
IBUF  _1775_ (
    .I(s15_data_i[19]),
    .O(_0146_[19])
  );
IBUF  _1776_ (
    .I(s15_data_i[2]),
    .O(_0146_[2])
  );
IBUF  _1777_ (
    .I(s15_data_i[20]),
    .O(_0146_[20])
  );
IBUF  _1778_ (
    .I(s15_data_i[21]),
    .O(_0146_[21])
  );
IBUF  _1779_ (
    .I(s15_data_i[22]),
    .O(_0146_[22])
  );
IBUF  _1780_ (
    .I(s15_data_i[23]),
    .O(_0146_[23])
  );
IBUF  _1781_ (
    .I(s15_data_i[24]),
    .O(_0146_[24])
  );
IBUF  _1782_ (
    .I(s15_data_i[25]),
    .O(_0146_[25])
  );
IBUF  _1783_ (
    .I(s15_data_i[26]),
    .O(_0146_[26])
  );
IBUF  _1784_ (
    .I(s15_data_i[27]),
    .O(_0146_[27])
  );
IBUF  _1785_ (
    .I(s15_data_i[28]),
    .O(_0146_[28])
  );
IBUF  _1786_ (
    .I(s15_data_i[29]),
    .O(_0146_[29])
  );
IBUF  _1787_ (
    .I(s15_data_i[3]),
    .O(_0146_[3])
  );
IBUF  _1788_ (
    .I(s15_data_i[30]),
    .O(_0146_[30])
  );
IBUF  _1789_ (
    .I(s15_data_i[31]),
    .O(_0146_[31])
  );
IBUF  _1790_ (
    .I(s15_data_i[4]),
    .O(_0146_[4])
  );
IBUF  _1791_ (
    .I(s15_data_i[5]),
    .O(_0146_[5])
  );
IBUF  _1792_ (
    .I(s15_data_i[6]),
    .O(_0146_[6])
  );
IBUF  _1793_ (
    .I(s15_data_i[7]),
    .O(_0146_[7])
  );
IBUF  _1794_ (
    .I(s15_data_i[8]),
    .O(_0146_[8])
  );
IBUF  _1795_ (
    .I(s15_data_i[9]),
    .O(_0146_[9])
  );
OBUF  _1796_ (
    .I(_0147_[0]),
    .O(s15_data_o[0])
  );
OBUF  _1797_ (
    .I(_0147_[1]),
    .O(s15_data_o[1])
  );
OBUF  _1798_ (
    .I(_0147_[10]),
    .O(s15_data_o[10])
  );
OBUF  _1799_ (
    .I(_0147_[11]),
    .O(s15_data_o[11])
  );
OBUF  _1800_ (
    .I(_0147_[12]),
    .O(s15_data_o[12])
  );
OBUF  _1801_ (
    .I(_0147_[13]),
    .O(s15_data_o[13])
  );
OBUF  _1802_ (
    .I(_0147_[14]),
    .O(s15_data_o[14])
  );
OBUF  _1803_ (
    .I(_0147_[15]),
    .O(s15_data_o[15])
  );
OBUF  _1804_ (
    .I(_0147_[16]),
    .O(s15_data_o[16])
  );
OBUF  _1805_ (
    .I(_0147_[17]),
    .O(s15_data_o[17])
  );
OBUF  _1806_ (
    .I(_0147_[18]),
    .O(s15_data_o[18])
  );
OBUF  _1807_ (
    .I(_0147_[19]),
    .O(s15_data_o[19])
  );
OBUF  _1808_ (
    .I(_0147_[2]),
    .O(s15_data_o[2])
  );
OBUF  _1809_ (
    .I(_0147_[20]),
    .O(s15_data_o[20])
  );
OBUF  _1810_ (
    .I(_0147_[21]),
    .O(s15_data_o[21])
  );
OBUF  _1811_ (
    .I(_0147_[22]),
    .O(s15_data_o[22])
  );
OBUF  _1812_ (
    .I(_0147_[23]),
    .O(s15_data_o[23])
  );
OBUF  _1813_ (
    .I(_0147_[24]),
    .O(s15_data_o[24])
  );
OBUF  _1814_ (
    .I(_0147_[25]),
    .O(s15_data_o[25])
  );
OBUF  _1815_ (
    .I(_0147_[26]),
    .O(s15_data_o[26])
  );
OBUF  _1816_ (
    .I(_0147_[27]),
    .O(s15_data_o[27])
  );
OBUF  _1817_ (
    .I(_0147_[28]),
    .O(s15_data_o[28])
  );
OBUF  _1818_ (
    .I(_0147_[29]),
    .O(s15_data_o[29])
  );
OBUF  _1819_ (
    .I(_0147_[3]),
    .O(s15_data_o[3])
  );
OBUF  _1820_ (
    .I(_0147_[30]),
    .O(s15_data_o[30])
  );
OBUF  _1821_ (
    .I(_0147_[31]),
    .O(s15_data_o[31])
  );
OBUF  _1822_ (
    .I(_0147_[4]),
    .O(s15_data_o[4])
  );
OBUF  _1823_ (
    .I(_0147_[5]),
    .O(s15_data_o[5])
  );
OBUF  _1824_ (
    .I(_0147_[6]),
    .O(s15_data_o[6])
  );
OBUF  _1825_ (
    .I(_0147_[7]),
    .O(s15_data_o[7])
  );
OBUF  _1826_ (
    .I(_0147_[8]),
    .O(s15_data_o[8])
  );
OBUF  _1827_ (
    .I(_0147_[9]),
    .O(s15_data_o[9])
  );
IBUF  _1828_ (
    .I(s15_err_i),
    .O(_0148_)
  );
IBUF  _1829_ (
    .I(s15_rty_i),
    .O(_0149_)
  );
OBUF  _1830_ (
    .I(_0150_[0]),
    .O(s15_sel_o[0])
  );
OBUF  _1831_ (
    .I(_0150_[1]),
    .O(s15_sel_o[1])
  );
OBUF  _1832_ (
    .I(_0150_[2]),
    .O(s15_sel_o[2])
  );
OBUF  _1833_ (
    .I(_0150_[3]),
    .O(s15_sel_o[3])
  );
OBUF  _1834_ (
    .I(_0151_),
    .O(s15_stb_o)
  );
OBUF  _1835_ (
    .I(_0152_),
    .O(s15_we_o)
  );
IBUF  _1836_ (
    .I(s1_ack_i),
    .O(_0153_)
  );
OBUF  _1837_ (
    .I(_0154_[0]),
    .O(s1_addr_o[0])
  );
OBUF  _1838_ (
    .I(_0154_[1]),
    .O(s1_addr_o[1])
  );
OBUF  _1839_ (
    .I(_0154_[10]),
    .O(s1_addr_o[10])
  );
OBUF  _1840_ (
    .I(_0154_[11]),
    .O(s1_addr_o[11])
  );
OBUF  _1841_ (
    .I(_0154_[12]),
    .O(s1_addr_o[12])
  );
OBUF  _1842_ (
    .I(_0154_[13]),
    .O(s1_addr_o[13])
  );
OBUF  _1843_ (
    .I(_0154_[14]),
    .O(s1_addr_o[14])
  );
OBUF  _1844_ (
    .I(_0154_[15]),
    .O(s1_addr_o[15])
  );
OBUF  _1845_ (
    .I(_0154_[16]),
    .O(s1_addr_o[16])
  );
OBUF  _1846_ (
    .I(_0154_[17]),
    .O(s1_addr_o[17])
  );
OBUF  _1847_ (
    .I(_0154_[18]),
    .O(s1_addr_o[18])
  );
OBUF  _1848_ (
    .I(_0154_[19]),
    .O(s1_addr_o[19])
  );
OBUF  _1849_ (
    .I(_0154_[2]),
    .O(s1_addr_o[2])
  );
OBUF  _1850_ (
    .I(_0154_[20]),
    .O(s1_addr_o[20])
  );
OBUF  _1851_ (
    .I(_0154_[21]),
    .O(s1_addr_o[21])
  );
OBUF  _1852_ (
    .I(_0154_[22]),
    .O(s1_addr_o[22])
  );
OBUF  _1853_ (
    .I(_0154_[23]),
    .O(s1_addr_o[23])
  );
OBUF  _1854_ (
    .I(_0154_[24]),
    .O(s1_addr_o[24])
  );
OBUF  _1855_ (
    .I(_0154_[25]),
    .O(s1_addr_o[25])
  );
OBUF  _1856_ (
    .I(_0154_[26]),
    .O(s1_addr_o[26])
  );
OBUF  _1857_ (
    .I(_0154_[27]),
    .O(s1_addr_o[27])
  );
OBUF  _1858_ (
    .I(_0154_[28]),
    .O(s1_addr_o[28])
  );
OBUF  _1859_ (
    .I(_0154_[29]),
    .O(s1_addr_o[29])
  );
OBUF  _1860_ (
    .I(_0154_[3]),
    .O(s1_addr_o[3])
  );
OBUF  _1861_ (
    .I(_0154_[30]),
    .O(s1_addr_o[30])
  );
OBUF  _1862_ (
    .I(_0154_[31]),
    .O(s1_addr_o[31])
  );
OBUF  _1863_ (
    .I(_0154_[4]),
    .O(s1_addr_o[4])
  );
OBUF  _1864_ (
    .I(_0154_[5]),
    .O(s1_addr_o[5])
  );
OBUF  _1865_ (
    .I(_0154_[6]),
    .O(s1_addr_o[6])
  );
OBUF  _1866_ (
    .I(_0154_[7]),
    .O(s1_addr_o[7])
  );
OBUF  _1867_ (
    .I(_0154_[8]),
    .O(s1_addr_o[8])
  );
OBUF  _1868_ (
    .I(_0154_[9]),
    .O(s1_addr_o[9])
  );
OBUF  _1869_ (
    .I(_0155_),
    .O(s1_cyc_o)
  );
IBUF  _1870_ (
    .I(s1_data_i[0]),
    .O(_0156_[0])
  );
IBUF  _1871_ (
    .I(s1_data_i[1]),
    .O(_0156_[1])
  );
IBUF  _1872_ (
    .I(s1_data_i[10]),
    .O(_0156_[10])
  );
IBUF  _1873_ (
    .I(s1_data_i[11]),
    .O(_0156_[11])
  );
IBUF  _1874_ (
    .I(s1_data_i[12]),
    .O(_0156_[12])
  );
IBUF  _1875_ (
    .I(s1_data_i[13]),
    .O(_0156_[13])
  );
IBUF  _1876_ (
    .I(s1_data_i[14]),
    .O(_0156_[14])
  );
IBUF  _1877_ (
    .I(s1_data_i[15]),
    .O(_0156_[15])
  );
IBUF  _1878_ (
    .I(s1_data_i[16]),
    .O(_0156_[16])
  );
IBUF  _1879_ (
    .I(s1_data_i[17]),
    .O(_0156_[17])
  );
IBUF  _1880_ (
    .I(s1_data_i[18]),
    .O(_0156_[18])
  );
IBUF  _1881_ (
    .I(s1_data_i[19]),
    .O(_0156_[19])
  );
IBUF  _1882_ (
    .I(s1_data_i[2]),
    .O(_0156_[2])
  );
IBUF  _1883_ (
    .I(s1_data_i[20]),
    .O(_0156_[20])
  );
IBUF  _1884_ (
    .I(s1_data_i[21]),
    .O(_0156_[21])
  );
IBUF  _1885_ (
    .I(s1_data_i[22]),
    .O(_0156_[22])
  );
IBUF  _1886_ (
    .I(s1_data_i[23]),
    .O(_0156_[23])
  );
IBUF  _1887_ (
    .I(s1_data_i[24]),
    .O(_0156_[24])
  );
IBUF  _1888_ (
    .I(s1_data_i[25]),
    .O(_0156_[25])
  );
IBUF  _1889_ (
    .I(s1_data_i[26]),
    .O(_0156_[26])
  );
IBUF  _1890_ (
    .I(s1_data_i[27]),
    .O(_0156_[27])
  );
IBUF  _1891_ (
    .I(s1_data_i[28]),
    .O(_0156_[28])
  );
IBUF  _1892_ (
    .I(s1_data_i[29]),
    .O(_0156_[29])
  );
IBUF  _1893_ (
    .I(s1_data_i[3]),
    .O(_0156_[3])
  );
IBUF  _1894_ (
    .I(s1_data_i[30]),
    .O(_0156_[30])
  );
IBUF  _1895_ (
    .I(s1_data_i[31]),
    .O(_0156_[31])
  );
IBUF  _1896_ (
    .I(s1_data_i[4]),
    .O(_0156_[4])
  );
IBUF  _1897_ (
    .I(s1_data_i[5]),
    .O(_0156_[5])
  );
IBUF  _1898_ (
    .I(s1_data_i[6]),
    .O(_0156_[6])
  );
IBUF  _1899_ (
    .I(s1_data_i[7]),
    .O(_0156_[7])
  );
IBUF  _1900_ (
    .I(s1_data_i[8]),
    .O(_0156_[8])
  );
IBUF  _1901_ (
    .I(s1_data_i[9]),
    .O(_0156_[9])
  );
OBUF  _1902_ (
    .I(_0157_[0]),
    .O(s1_data_o[0])
  );
OBUF  _1903_ (
    .I(_0157_[1]),
    .O(s1_data_o[1])
  );
OBUF  _1904_ (
    .I(_0157_[10]),
    .O(s1_data_o[10])
  );
OBUF  _1905_ (
    .I(_0157_[11]),
    .O(s1_data_o[11])
  );
OBUF  _1906_ (
    .I(_0157_[12]),
    .O(s1_data_o[12])
  );
OBUF  _1907_ (
    .I(_0157_[13]),
    .O(s1_data_o[13])
  );
OBUF  _1908_ (
    .I(_0157_[14]),
    .O(s1_data_o[14])
  );
OBUF  _1909_ (
    .I(_0157_[15]),
    .O(s1_data_o[15])
  );
OBUF  _1910_ (
    .I(_0157_[16]),
    .O(s1_data_o[16])
  );
OBUF  _1911_ (
    .I(_0157_[17]),
    .O(s1_data_o[17])
  );
OBUF  _1912_ (
    .I(_0157_[18]),
    .O(s1_data_o[18])
  );
OBUF  _1913_ (
    .I(_0157_[19]),
    .O(s1_data_o[19])
  );
OBUF  _1914_ (
    .I(_0157_[2]),
    .O(s1_data_o[2])
  );
OBUF  _1915_ (
    .I(_0157_[20]),
    .O(s1_data_o[20])
  );
OBUF  _1916_ (
    .I(_0157_[21]),
    .O(s1_data_o[21])
  );
OBUF  _1917_ (
    .I(_0157_[22]),
    .O(s1_data_o[22])
  );
OBUF  _1918_ (
    .I(_0157_[23]),
    .O(s1_data_o[23])
  );
OBUF  _1919_ (
    .I(_0157_[24]),
    .O(s1_data_o[24])
  );
OBUF  _1920_ (
    .I(_0157_[25]),
    .O(s1_data_o[25])
  );
OBUF  _1921_ (
    .I(_0157_[26]),
    .O(s1_data_o[26])
  );
OBUF  _1922_ (
    .I(_0157_[27]),
    .O(s1_data_o[27])
  );
OBUF  _1923_ (
    .I(_0157_[28]),
    .O(s1_data_o[28])
  );
OBUF  _1924_ (
    .I(_0157_[29]),
    .O(s1_data_o[29])
  );
OBUF  _1925_ (
    .I(_0157_[3]),
    .O(s1_data_o[3])
  );
OBUF  _1926_ (
    .I(_0157_[30]),
    .O(s1_data_o[30])
  );
OBUF  _1927_ (
    .I(_0157_[31]),
    .O(s1_data_o[31])
  );
OBUF  _1928_ (
    .I(_0157_[4]),
    .O(s1_data_o[4])
  );
OBUF  _1929_ (
    .I(_0157_[5]),
    .O(s1_data_o[5])
  );
OBUF  _1930_ (
    .I(_0157_[6]),
    .O(s1_data_o[6])
  );
OBUF  _1931_ (
    .I(_0157_[7]),
    .O(s1_data_o[7])
  );
OBUF  _1932_ (
    .I(_0157_[8]),
    .O(s1_data_o[8])
  );
OBUF  _1933_ (
    .I(_0157_[9]),
    .O(s1_data_o[9])
  );
IBUF  _1934_ (
    .I(s1_err_i),
    .O(_0158_)
  );
IBUF  _1935_ (
    .I(s1_rty_i),
    .O(_0159_)
  );
OBUF  _1936_ (
    .I(_0160_[0]),
    .O(s1_sel_o[0])
  );
OBUF  _1937_ (
    .I(_0160_[1]),
    .O(s1_sel_o[1])
  );
OBUF  _1938_ (
    .I(_0160_[2]),
    .O(s1_sel_o[2])
  );
OBUF  _1939_ (
    .I(_0160_[3]),
    .O(s1_sel_o[3])
  );
OBUF  _1940_ (
    .I(_0161_),
    .O(s1_stb_o)
  );
OBUF  _1941_ (
    .I(_0162_),
    .O(s1_we_o)
  );
IBUF  _1942_ (
    .I(s2_ack_i),
    .O(_0163_)
  );
OBUF  _1943_ (
    .I(_0164_[0]),
    .O(s2_addr_o[0])
  );
OBUF  _1944_ (
    .I(_0164_[1]),
    .O(s2_addr_o[1])
  );
OBUF  _1945_ (
    .I(_0164_[10]),
    .O(s2_addr_o[10])
  );
OBUF  _1946_ (
    .I(_0164_[11]),
    .O(s2_addr_o[11])
  );
OBUF  _1947_ (
    .I(_0164_[12]),
    .O(s2_addr_o[12])
  );
OBUF  _1948_ (
    .I(_0164_[13]),
    .O(s2_addr_o[13])
  );
OBUF  _1949_ (
    .I(_0164_[14]),
    .O(s2_addr_o[14])
  );
OBUF  _1950_ (
    .I(_0164_[15]),
    .O(s2_addr_o[15])
  );
OBUF  _1951_ (
    .I(_0164_[16]),
    .O(s2_addr_o[16])
  );
OBUF  _1952_ (
    .I(_0164_[17]),
    .O(s2_addr_o[17])
  );
OBUF  _1953_ (
    .I(_0164_[18]),
    .O(s2_addr_o[18])
  );
OBUF  _1954_ (
    .I(_0164_[19]),
    .O(s2_addr_o[19])
  );
OBUF  _1955_ (
    .I(_0164_[2]),
    .O(s2_addr_o[2])
  );
OBUF  _1956_ (
    .I(_0164_[20]),
    .O(s2_addr_o[20])
  );
OBUF  _1957_ (
    .I(_0164_[21]),
    .O(s2_addr_o[21])
  );
OBUF  _1958_ (
    .I(_0164_[22]),
    .O(s2_addr_o[22])
  );
OBUF  _1959_ (
    .I(_0164_[23]),
    .O(s2_addr_o[23])
  );
OBUF  _1960_ (
    .I(_0164_[24]),
    .O(s2_addr_o[24])
  );
OBUF  _1961_ (
    .I(_0164_[25]),
    .O(s2_addr_o[25])
  );
OBUF  _1962_ (
    .I(_0164_[26]),
    .O(s2_addr_o[26])
  );
OBUF  _1963_ (
    .I(_0164_[27]),
    .O(s2_addr_o[27])
  );
OBUF  _1964_ (
    .I(_0164_[28]),
    .O(s2_addr_o[28])
  );
OBUF  _1965_ (
    .I(_0164_[29]),
    .O(s2_addr_o[29])
  );
OBUF  _1966_ (
    .I(_0164_[3]),
    .O(s2_addr_o[3])
  );
OBUF  _1967_ (
    .I(_0164_[30]),
    .O(s2_addr_o[30])
  );
OBUF  _1968_ (
    .I(_0164_[31]),
    .O(s2_addr_o[31])
  );
OBUF  _1969_ (
    .I(_0164_[4]),
    .O(s2_addr_o[4])
  );
OBUF  _1970_ (
    .I(_0164_[5]),
    .O(s2_addr_o[5])
  );
OBUF  _1971_ (
    .I(_0164_[6]),
    .O(s2_addr_o[6])
  );
OBUF  _1972_ (
    .I(_0164_[7]),
    .O(s2_addr_o[7])
  );
OBUF  _1973_ (
    .I(_0164_[8]),
    .O(s2_addr_o[8])
  );
OBUF  _1974_ (
    .I(_0164_[9]),
    .O(s2_addr_o[9])
  );
OBUF  _1975_ (
    .I(_0165_),
    .O(s2_cyc_o)
  );
IBUF  _1976_ (
    .I(s2_data_i[0]),
    .O(_0166_[0])
  );
IBUF  _1977_ (
    .I(s2_data_i[1]),
    .O(_0166_[1])
  );
IBUF  _1978_ (
    .I(s2_data_i[10]),
    .O(_0166_[10])
  );
IBUF  _1979_ (
    .I(s2_data_i[11]),
    .O(_0166_[11])
  );
IBUF  _1980_ (
    .I(s2_data_i[12]),
    .O(_0166_[12])
  );
IBUF  _1981_ (
    .I(s2_data_i[13]),
    .O(_0166_[13])
  );
IBUF  _1982_ (
    .I(s2_data_i[14]),
    .O(_0166_[14])
  );
IBUF  _1983_ (
    .I(s2_data_i[15]),
    .O(_0166_[15])
  );
IBUF  _1984_ (
    .I(s2_data_i[16]),
    .O(_0166_[16])
  );
IBUF  _1985_ (
    .I(s2_data_i[17]),
    .O(_0166_[17])
  );
IBUF  _1986_ (
    .I(s2_data_i[18]),
    .O(_0166_[18])
  );
IBUF  _1987_ (
    .I(s2_data_i[19]),
    .O(_0166_[19])
  );
IBUF  _1988_ (
    .I(s2_data_i[2]),
    .O(_0166_[2])
  );
IBUF  _1989_ (
    .I(s2_data_i[20]),
    .O(_0166_[20])
  );
IBUF  _1990_ (
    .I(s2_data_i[21]),
    .O(_0166_[21])
  );
IBUF  _1991_ (
    .I(s2_data_i[22]),
    .O(_0166_[22])
  );
IBUF  _1992_ (
    .I(s2_data_i[23]),
    .O(_0166_[23])
  );
IBUF  _1993_ (
    .I(s2_data_i[24]),
    .O(_0166_[24])
  );
IBUF  _1994_ (
    .I(s2_data_i[25]),
    .O(_0166_[25])
  );
IBUF  _1995_ (
    .I(s2_data_i[26]),
    .O(_0166_[26])
  );
IBUF  _1996_ (
    .I(s2_data_i[27]),
    .O(_0166_[27])
  );
IBUF  _1997_ (
    .I(s2_data_i[28]),
    .O(_0166_[28])
  );
IBUF  _1998_ (
    .I(s2_data_i[29]),
    .O(_0166_[29])
  );
IBUF  _1999_ (
    .I(s2_data_i[3]),
    .O(_0166_[3])
  );
IBUF  _2000_ (
    .I(s2_data_i[30]),
    .O(_0166_[30])
  );
IBUF  _2001_ (
    .I(s2_data_i[31]),
    .O(_0166_[31])
  );
IBUF  _2002_ (
    .I(s2_data_i[4]),
    .O(_0166_[4])
  );
IBUF  _2003_ (
    .I(s2_data_i[5]),
    .O(_0166_[5])
  );
IBUF  _2004_ (
    .I(s2_data_i[6]),
    .O(_0166_[6])
  );
IBUF  _2005_ (
    .I(s2_data_i[7]),
    .O(_0166_[7])
  );
IBUF  _2006_ (
    .I(s2_data_i[8]),
    .O(_0166_[8])
  );
IBUF  _2007_ (
    .I(s2_data_i[9]),
    .O(_0166_[9])
  );
OBUF  _2008_ (
    .I(_0167_[0]),
    .O(s2_data_o[0])
  );
OBUF  _2009_ (
    .I(_0167_[1]),
    .O(s2_data_o[1])
  );
OBUF  _2010_ (
    .I(_0167_[10]),
    .O(s2_data_o[10])
  );
OBUF  _2011_ (
    .I(_0167_[11]),
    .O(s2_data_o[11])
  );
OBUF  _2012_ (
    .I(_0167_[12]),
    .O(s2_data_o[12])
  );
OBUF  _2013_ (
    .I(_0167_[13]),
    .O(s2_data_o[13])
  );
OBUF  _2014_ (
    .I(_0167_[14]),
    .O(s2_data_o[14])
  );
OBUF  _2015_ (
    .I(_0167_[15]),
    .O(s2_data_o[15])
  );
OBUF  _2016_ (
    .I(_0167_[16]),
    .O(s2_data_o[16])
  );
OBUF  _2017_ (
    .I(_0167_[17]),
    .O(s2_data_o[17])
  );
OBUF  _2018_ (
    .I(_0167_[18]),
    .O(s2_data_o[18])
  );
OBUF  _2019_ (
    .I(_0167_[19]),
    .O(s2_data_o[19])
  );
OBUF  _2020_ (
    .I(_0167_[2]),
    .O(s2_data_o[2])
  );
OBUF  _2021_ (
    .I(_0167_[20]),
    .O(s2_data_o[20])
  );
OBUF  _2022_ (
    .I(_0167_[21]),
    .O(s2_data_o[21])
  );
OBUF  _2023_ (
    .I(_0167_[22]),
    .O(s2_data_o[22])
  );
OBUF  _2024_ (
    .I(_0167_[23]),
    .O(s2_data_o[23])
  );
OBUF  _2025_ (
    .I(_0167_[24]),
    .O(s2_data_o[24])
  );
OBUF  _2026_ (
    .I(_0167_[25]),
    .O(s2_data_o[25])
  );
OBUF  _2027_ (
    .I(_0167_[26]),
    .O(s2_data_o[26])
  );
OBUF  _2028_ (
    .I(_0167_[27]),
    .O(s2_data_o[27])
  );
OBUF  _2029_ (
    .I(_0167_[28]),
    .O(s2_data_o[28])
  );
OBUF  _2030_ (
    .I(_0167_[29]),
    .O(s2_data_o[29])
  );
OBUF  _2031_ (
    .I(_0167_[3]),
    .O(s2_data_o[3])
  );
OBUF  _2032_ (
    .I(_0167_[30]),
    .O(s2_data_o[30])
  );
OBUF  _2033_ (
    .I(_0167_[31]),
    .O(s2_data_o[31])
  );
OBUF  _2034_ (
    .I(_0167_[4]),
    .O(s2_data_o[4])
  );
OBUF  _2035_ (
    .I(_0167_[5]),
    .O(s2_data_o[5])
  );
OBUF  _2036_ (
    .I(_0167_[6]),
    .O(s2_data_o[6])
  );
OBUF  _2037_ (
    .I(_0167_[7]),
    .O(s2_data_o[7])
  );
OBUF  _2038_ (
    .I(_0167_[8]),
    .O(s2_data_o[8])
  );
OBUF  _2039_ (
    .I(_0167_[9]),
    .O(s2_data_o[9])
  );
IBUF  _2040_ (
    .I(s2_err_i),
    .O(_0168_)
  );
IBUF  _2041_ (
    .I(s2_rty_i),
    .O(_0169_)
  );
OBUF  _2042_ (
    .I(_0170_[0]),
    .O(s2_sel_o[0])
  );
OBUF  _2043_ (
    .I(_0170_[1]),
    .O(s2_sel_o[1])
  );
OBUF  _2044_ (
    .I(_0170_[2]),
    .O(s2_sel_o[2])
  );
OBUF  _2045_ (
    .I(_0170_[3]),
    .O(s2_sel_o[3])
  );
OBUF  _2046_ (
    .I(_0171_),
    .O(s2_stb_o)
  );
OBUF  _2047_ (
    .I(_0172_),
    .O(s2_we_o)
  );
IBUF  _2048_ (
    .I(s3_ack_i),
    .O(_0173_)
  );
OBUF  _2049_ (
    .I(_0174_[0]),
    .O(s3_addr_o[0])
  );
OBUF  _2050_ (
    .I(_0174_[1]),
    .O(s3_addr_o[1])
  );
OBUF  _2051_ (
    .I(_0174_[10]),
    .O(s3_addr_o[10])
  );
OBUF  _2052_ (
    .I(_0174_[11]),
    .O(s3_addr_o[11])
  );
OBUF  _2053_ (
    .I(_0174_[12]),
    .O(s3_addr_o[12])
  );
OBUF  _2054_ (
    .I(_0174_[13]),
    .O(s3_addr_o[13])
  );
OBUF  _2055_ (
    .I(_0174_[14]),
    .O(s3_addr_o[14])
  );
OBUF  _2056_ (
    .I(_0174_[15]),
    .O(s3_addr_o[15])
  );
OBUF  _2057_ (
    .I(_0174_[16]),
    .O(s3_addr_o[16])
  );
OBUF  _2058_ (
    .I(_0174_[17]),
    .O(s3_addr_o[17])
  );
OBUF  _2059_ (
    .I(_0174_[18]),
    .O(s3_addr_o[18])
  );
OBUF  _2060_ (
    .I(_0174_[19]),
    .O(s3_addr_o[19])
  );
OBUF  _2061_ (
    .I(_0174_[2]),
    .O(s3_addr_o[2])
  );
OBUF  _2062_ (
    .I(_0174_[20]),
    .O(s3_addr_o[20])
  );
OBUF  _2063_ (
    .I(_0174_[21]),
    .O(s3_addr_o[21])
  );
OBUF  _2064_ (
    .I(_0174_[22]),
    .O(s3_addr_o[22])
  );
OBUF  _2065_ (
    .I(_0174_[23]),
    .O(s3_addr_o[23])
  );
OBUF  _2066_ (
    .I(_0174_[24]),
    .O(s3_addr_o[24])
  );
OBUF  _2067_ (
    .I(_0174_[25]),
    .O(s3_addr_o[25])
  );
OBUF  _2068_ (
    .I(_0174_[26]),
    .O(s3_addr_o[26])
  );
OBUF  _2069_ (
    .I(_0174_[27]),
    .O(s3_addr_o[27])
  );
OBUF  _2070_ (
    .I(_0174_[28]),
    .O(s3_addr_o[28])
  );
OBUF  _2071_ (
    .I(_0174_[29]),
    .O(s3_addr_o[29])
  );
OBUF  _2072_ (
    .I(_0174_[3]),
    .O(s3_addr_o[3])
  );
OBUF  _2073_ (
    .I(_0174_[30]),
    .O(s3_addr_o[30])
  );
OBUF  _2074_ (
    .I(_0174_[31]),
    .O(s3_addr_o[31])
  );
OBUF  _2075_ (
    .I(_0174_[4]),
    .O(s3_addr_o[4])
  );
OBUF  _2076_ (
    .I(_0174_[5]),
    .O(s3_addr_o[5])
  );
OBUF  _2077_ (
    .I(_0174_[6]),
    .O(s3_addr_o[6])
  );
OBUF  _2078_ (
    .I(_0174_[7]),
    .O(s3_addr_o[7])
  );
OBUF  _2079_ (
    .I(_0174_[8]),
    .O(s3_addr_o[8])
  );
OBUF  _2080_ (
    .I(_0174_[9]),
    .O(s3_addr_o[9])
  );
OBUF  _2081_ (
    .I(_0175_),
    .O(s3_cyc_o)
  );
IBUF  _2082_ (
    .I(s3_data_i[0]),
    .O(_0176_[0])
  );
IBUF  _2083_ (
    .I(s3_data_i[1]),
    .O(_0176_[1])
  );
IBUF  _2084_ (
    .I(s3_data_i[10]),
    .O(_0176_[10])
  );
IBUF  _2085_ (
    .I(s3_data_i[11]),
    .O(_0176_[11])
  );
IBUF  _2086_ (
    .I(s3_data_i[12]),
    .O(_0176_[12])
  );
IBUF  _2087_ (
    .I(s3_data_i[13]),
    .O(_0176_[13])
  );
IBUF  _2088_ (
    .I(s3_data_i[14]),
    .O(_0176_[14])
  );
IBUF  _2089_ (
    .I(s3_data_i[15]),
    .O(_0176_[15])
  );
IBUF  _2090_ (
    .I(s3_data_i[16]),
    .O(_0176_[16])
  );
IBUF  _2091_ (
    .I(s3_data_i[17]),
    .O(_0176_[17])
  );
IBUF  _2092_ (
    .I(s3_data_i[18]),
    .O(_0176_[18])
  );
IBUF  _2093_ (
    .I(s3_data_i[19]),
    .O(_0176_[19])
  );
IBUF  _2094_ (
    .I(s3_data_i[2]),
    .O(_0176_[2])
  );
IBUF  _2095_ (
    .I(s3_data_i[20]),
    .O(_0176_[20])
  );
IBUF  _2096_ (
    .I(s3_data_i[21]),
    .O(_0176_[21])
  );
IBUF  _2097_ (
    .I(s3_data_i[22]),
    .O(_0176_[22])
  );
IBUF  _2098_ (
    .I(s3_data_i[23]),
    .O(_0176_[23])
  );
IBUF  _2099_ (
    .I(s3_data_i[24]),
    .O(_0176_[24])
  );
IBUF  _2100_ (
    .I(s3_data_i[25]),
    .O(_0176_[25])
  );
IBUF  _2101_ (
    .I(s3_data_i[26]),
    .O(_0176_[26])
  );
IBUF  _2102_ (
    .I(s3_data_i[27]),
    .O(_0176_[27])
  );
IBUF  _2103_ (
    .I(s3_data_i[28]),
    .O(_0176_[28])
  );
IBUF  _2104_ (
    .I(s3_data_i[29]),
    .O(_0176_[29])
  );
IBUF  _2105_ (
    .I(s3_data_i[3]),
    .O(_0176_[3])
  );
IBUF  _2106_ (
    .I(s3_data_i[30]),
    .O(_0176_[30])
  );
IBUF  _2107_ (
    .I(s3_data_i[31]),
    .O(_0176_[31])
  );
IBUF  _2108_ (
    .I(s3_data_i[4]),
    .O(_0176_[4])
  );
IBUF  _2109_ (
    .I(s3_data_i[5]),
    .O(_0176_[5])
  );
IBUF  _2110_ (
    .I(s3_data_i[6]),
    .O(_0176_[6])
  );
IBUF  _2111_ (
    .I(s3_data_i[7]),
    .O(_0176_[7])
  );
IBUF  _2112_ (
    .I(s3_data_i[8]),
    .O(_0176_[8])
  );
IBUF  _2113_ (
    .I(s3_data_i[9]),
    .O(_0176_[9])
  );
OBUF  _2114_ (
    .I(_0177_[0]),
    .O(s3_data_o[0])
  );
OBUF  _2115_ (
    .I(_0177_[1]),
    .O(s3_data_o[1])
  );
OBUF  _2116_ (
    .I(_0177_[10]),
    .O(s3_data_o[10])
  );
OBUF  _2117_ (
    .I(_0177_[11]),
    .O(s3_data_o[11])
  );
OBUF  _2118_ (
    .I(_0177_[12]),
    .O(s3_data_o[12])
  );
OBUF  _2119_ (
    .I(_0177_[13]),
    .O(s3_data_o[13])
  );
OBUF  _2120_ (
    .I(_0177_[14]),
    .O(s3_data_o[14])
  );
OBUF  _2121_ (
    .I(_0177_[15]),
    .O(s3_data_o[15])
  );
OBUF  _2122_ (
    .I(_0177_[16]),
    .O(s3_data_o[16])
  );
OBUF  _2123_ (
    .I(_0177_[17]),
    .O(s3_data_o[17])
  );
OBUF  _2124_ (
    .I(_0177_[18]),
    .O(s3_data_o[18])
  );
OBUF  _2125_ (
    .I(_0177_[19]),
    .O(s3_data_o[19])
  );
OBUF  _2126_ (
    .I(_0177_[2]),
    .O(s3_data_o[2])
  );
OBUF  _2127_ (
    .I(_0177_[20]),
    .O(s3_data_o[20])
  );
OBUF  _2128_ (
    .I(_0177_[21]),
    .O(s3_data_o[21])
  );
OBUF  _2129_ (
    .I(_0177_[22]),
    .O(s3_data_o[22])
  );
OBUF  _2130_ (
    .I(_0177_[23]),
    .O(s3_data_o[23])
  );
OBUF  _2131_ (
    .I(_0177_[24]),
    .O(s3_data_o[24])
  );
OBUF  _2132_ (
    .I(_0177_[25]),
    .O(s3_data_o[25])
  );
OBUF  _2133_ (
    .I(_0177_[26]),
    .O(s3_data_o[26])
  );
OBUF  _2134_ (
    .I(_0177_[27]),
    .O(s3_data_o[27])
  );
OBUF  _2135_ (
    .I(_0177_[28]),
    .O(s3_data_o[28])
  );
OBUF  _2136_ (
    .I(_0177_[29]),
    .O(s3_data_o[29])
  );
OBUF  _2137_ (
    .I(_0177_[3]),
    .O(s3_data_o[3])
  );
OBUF  _2138_ (
    .I(_0177_[30]),
    .O(s3_data_o[30])
  );
OBUF  _2139_ (
    .I(_0177_[31]),
    .O(s3_data_o[31])
  );
OBUF  _2140_ (
    .I(_0177_[4]),
    .O(s3_data_o[4])
  );
OBUF  _2141_ (
    .I(_0177_[5]),
    .O(s3_data_o[5])
  );
OBUF  _2142_ (
    .I(_0177_[6]),
    .O(s3_data_o[6])
  );
OBUF  _2143_ (
    .I(_0177_[7]),
    .O(s3_data_o[7])
  );
OBUF  _2144_ (
    .I(_0177_[8]),
    .O(s3_data_o[8])
  );
OBUF  _2145_ (
    .I(_0177_[9]),
    .O(s3_data_o[9])
  );
IBUF  _2146_ (
    .I(s3_err_i),
    .O(_0178_)
  );
IBUF  _2147_ (
    .I(s3_rty_i),
    .O(_0179_)
  );
OBUF  _2148_ (
    .I(_0180_[0]),
    .O(s3_sel_o[0])
  );
OBUF  _2149_ (
    .I(_0180_[1]),
    .O(s3_sel_o[1])
  );
OBUF  _2150_ (
    .I(_0180_[2]),
    .O(s3_sel_o[2])
  );
OBUF  _2151_ (
    .I(_0180_[3]),
    .O(s3_sel_o[3])
  );
OBUF  _2152_ (
    .I(_0181_),
    .O(s3_stb_o)
  );
OBUF  _2153_ (
    .I(_0182_),
    .O(s3_we_o)
  );
IBUF  _2154_ (
    .I(s4_ack_i),
    .O(_0183_)
  );
OBUF  _2155_ (
    .I(_0184_[0]),
    .O(s4_addr_o[0])
  );
OBUF  _2156_ (
    .I(_0184_[1]),
    .O(s4_addr_o[1])
  );
OBUF  _2157_ (
    .I(_0184_[10]),
    .O(s4_addr_o[10])
  );
OBUF  _2158_ (
    .I(_0184_[11]),
    .O(s4_addr_o[11])
  );
OBUF  _2159_ (
    .I(_0184_[12]),
    .O(s4_addr_o[12])
  );
OBUF  _2160_ (
    .I(_0184_[13]),
    .O(s4_addr_o[13])
  );
OBUF  _2161_ (
    .I(_0184_[14]),
    .O(s4_addr_o[14])
  );
OBUF  _2162_ (
    .I(_0184_[15]),
    .O(s4_addr_o[15])
  );
OBUF  _2163_ (
    .I(_0184_[16]),
    .O(s4_addr_o[16])
  );
OBUF  _2164_ (
    .I(_0184_[17]),
    .O(s4_addr_o[17])
  );
OBUF  _2165_ (
    .I(_0184_[18]),
    .O(s4_addr_o[18])
  );
OBUF  _2166_ (
    .I(_0184_[19]),
    .O(s4_addr_o[19])
  );
OBUF  _2167_ (
    .I(_0184_[2]),
    .O(s4_addr_o[2])
  );
OBUF  _2168_ (
    .I(_0184_[20]),
    .O(s4_addr_o[20])
  );
OBUF  _2169_ (
    .I(_0184_[21]),
    .O(s4_addr_o[21])
  );
OBUF  _2170_ (
    .I(_0184_[22]),
    .O(s4_addr_o[22])
  );
OBUF  _2171_ (
    .I(_0184_[23]),
    .O(s4_addr_o[23])
  );
OBUF  _2172_ (
    .I(_0184_[24]),
    .O(s4_addr_o[24])
  );
OBUF  _2173_ (
    .I(_0184_[25]),
    .O(s4_addr_o[25])
  );
OBUF  _2174_ (
    .I(_0184_[26]),
    .O(s4_addr_o[26])
  );
OBUF  _2175_ (
    .I(_0184_[27]),
    .O(s4_addr_o[27])
  );
OBUF  _2176_ (
    .I(_0184_[28]),
    .O(s4_addr_o[28])
  );
OBUF  _2177_ (
    .I(_0184_[29]),
    .O(s4_addr_o[29])
  );
OBUF  _2178_ (
    .I(_0184_[3]),
    .O(s4_addr_o[3])
  );
OBUF  _2179_ (
    .I(_0184_[30]),
    .O(s4_addr_o[30])
  );
OBUF  _2180_ (
    .I(_0184_[31]),
    .O(s4_addr_o[31])
  );
OBUF  _2181_ (
    .I(_0184_[4]),
    .O(s4_addr_o[4])
  );
OBUF  _2182_ (
    .I(_0184_[5]),
    .O(s4_addr_o[5])
  );
OBUF  _2183_ (
    .I(_0184_[6]),
    .O(s4_addr_o[6])
  );
OBUF  _2184_ (
    .I(_0184_[7]),
    .O(s4_addr_o[7])
  );
OBUF  _2185_ (
    .I(_0184_[8]),
    .O(s4_addr_o[8])
  );
OBUF  _2186_ (
    .I(_0184_[9]),
    .O(s4_addr_o[9])
  );
OBUF  _2187_ (
    .I(_0185_),
    .O(s4_cyc_o)
  );
IBUF  _2188_ (
    .I(s4_data_i[0]),
    .O(_0186_[0])
  );
IBUF  _2189_ (
    .I(s4_data_i[1]),
    .O(_0186_[1])
  );
IBUF  _2190_ (
    .I(s4_data_i[10]),
    .O(_0186_[10])
  );
IBUF  _2191_ (
    .I(s4_data_i[11]),
    .O(_0186_[11])
  );
IBUF  _2192_ (
    .I(s4_data_i[12]),
    .O(_0186_[12])
  );
IBUF  _2193_ (
    .I(s4_data_i[13]),
    .O(_0186_[13])
  );
IBUF  _2194_ (
    .I(s4_data_i[14]),
    .O(_0186_[14])
  );
IBUF  _2195_ (
    .I(s4_data_i[15]),
    .O(_0186_[15])
  );
IBUF  _2196_ (
    .I(s4_data_i[16]),
    .O(_0186_[16])
  );
IBUF  _2197_ (
    .I(s4_data_i[17]),
    .O(_0186_[17])
  );
IBUF  _2198_ (
    .I(s4_data_i[18]),
    .O(_0186_[18])
  );
IBUF  _2199_ (
    .I(s4_data_i[19]),
    .O(_0186_[19])
  );
IBUF  _2200_ (
    .I(s4_data_i[2]),
    .O(_0186_[2])
  );
IBUF  _2201_ (
    .I(s4_data_i[20]),
    .O(_0186_[20])
  );
IBUF  _2202_ (
    .I(s4_data_i[21]),
    .O(_0186_[21])
  );
IBUF  _2203_ (
    .I(s4_data_i[22]),
    .O(_0186_[22])
  );
IBUF  _2204_ (
    .I(s4_data_i[23]),
    .O(_0186_[23])
  );
IBUF  _2205_ (
    .I(s4_data_i[24]),
    .O(_0186_[24])
  );
IBUF  _2206_ (
    .I(s4_data_i[25]),
    .O(_0186_[25])
  );
IBUF  _2207_ (
    .I(s4_data_i[26]),
    .O(_0186_[26])
  );
IBUF  _2208_ (
    .I(s4_data_i[27]),
    .O(_0186_[27])
  );
IBUF  _2209_ (
    .I(s4_data_i[28]),
    .O(_0186_[28])
  );
IBUF  _2210_ (
    .I(s4_data_i[29]),
    .O(_0186_[29])
  );
IBUF  _2211_ (
    .I(s4_data_i[3]),
    .O(_0186_[3])
  );
IBUF  _2212_ (
    .I(s4_data_i[30]),
    .O(_0186_[30])
  );
IBUF  _2213_ (
    .I(s4_data_i[31]),
    .O(_0186_[31])
  );
IBUF  _2214_ (
    .I(s4_data_i[4]),
    .O(_0186_[4])
  );
IBUF  _2215_ (
    .I(s4_data_i[5]),
    .O(_0186_[5])
  );
IBUF  _2216_ (
    .I(s4_data_i[6]),
    .O(_0186_[6])
  );
IBUF  _2217_ (
    .I(s4_data_i[7]),
    .O(_0186_[7])
  );
IBUF  _2218_ (
    .I(s4_data_i[8]),
    .O(_0186_[8])
  );
IBUF  _2219_ (
    .I(s4_data_i[9]),
    .O(_0186_[9])
  );
OBUF  _2220_ (
    .I(_0187_[0]),
    .O(s4_data_o[0])
  );
OBUF  _2221_ (
    .I(_0187_[1]),
    .O(s4_data_o[1])
  );
OBUF  _2222_ (
    .I(_0187_[10]),
    .O(s4_data_o[10])
  );
OBUF  _2223_ (
    .I(_0187_[11]),
    .O(s4_data_o[11])
  );
OBUF  _2224_ (
    .I(_0187_[12]),
    .O(s4_data_o[12])
  );
OBUF  _2225_ (
    .I(_0187_[13]),
    .O(s4_data_o[13])
  );
OBUF  _2226_ (
    .I(_0187_[14]),
    .O(s4_data_o[14])
  );
OBUF  _2227_ (
    .I(_0187_[15]),
    .O(s4_data_o[15])
  );
OBUF  _2228_ (
    .I(_0187_[16]),
    .O(s4_data_o[16])
  );
OBUF  _2229_ (
    .I(_0187_[17]),
    .O(s4_data_o[17])
  );
OBUF  _2230_ (
    .I(_0187_[18]),
    .O(s4_data_o[18])
  );
OBUF  _2231_ (
    .I(_0187_[19]),
    .O(s4_data_o[19])
  );
OBUF  _2232_ (
    .I(_0187_[2]),
    .O(s4_data_o[2])
  );
OBUF  _2233_ (
    .I(_0187_[20]),
    .O(s4_data_o[20])
  );
OBUF  _2234_ (
    .I(_0187_[21]),
    .O(s4_data_o[21])
  );
OBUF  _2235_ (
    .I(_0187_[22]),
    .O(s4_data_o[22])
  );
OBUF  _2236_ (
    .I(_0187_[23]),
    .O(s4_data_o[23])
  );
OBUF  _2237_ (
    .I(_0187_[24]),
    .O(s4_data_o[24])
  );
OBUF  _2238_ (
    .I(_0187_[25]),
    .O(s4_data_o[25])
  );
OBUF  _2239_ (
    .I(_0187_[26]),
    .O(s4_data_o[26])
  );
OBUF  _2240_ (
    .I(_0187_[27]),
    .O(s4_data_o[27])
  );
OBUF  _2241_ (
    .I(_0187_[28]),
    .O(s4_data_o[28])
  );
OBUF  _2242_ (
    .I(_0187_[29]),
    .O(s4_data_o[29])
  );
OBUF  _2243_ (
    .I(_0187_[3]),
    .O(s4_data_o[3])
  );
OBUF  _2244_ (
    .I(_0187_[30]),
    .O(s4_data_o[30])
  );
OBUF  _2245_ (
    .I(_0187_[31]),
    .O(s4_data_o[31])
  );
OBUF  _2246_ (
    .I(_0187_[4]),
    .O(s4_data_o[4])
  );
OBUF  _2247_ (
    .I(_0187_[5]),
    .O(s4_data_o[5])
  );
OBUF  _2248_ (
    .I(_0187_[6]),
    .O(s4_data_o[6])
  );
OBUF  _2249_ (
    .I(_0187_[7]),
    .O(s4_data_o[7])
  );
OBUF  _2250_ (
    .I(_0187_[8]),
    .O(s4_data_o[8])
  );
OBUF  _2251_ (
    .I(_0187_[9]),
    .O(s4_data_o[9])
  );
IBUF  _2252_ (
    .I(s4_err_i),
    .O(_0188_)
  );
IBUF  _2253_ (
    .I(s4_rty_i),
    .O(_0189_)
  );
OBUF  _2254_ (
    .I(_0190_[0]),
    .O(s4_sel_o[0])
  );
OBUF  _2255_ (
    .I(_0190_[1]),
    .O(s4_sel_o[1])
  );
OBUF  _2256_ (
    .I(_0190_[2]),
    .O(s4_sel_o[2])
  );
OBUF  _2257_ (
    .I(_0190_[3]),
    .O(s4_sel_o[3])
  );
OBUF  _2258_ (
    .I(_0191_),
    .O(s4_stb_o)
  );
OBUF  _2259_ (
    .I(_0192_),
    .O(s4_we_o)
  );
IBUF  _2260_ (
    .I(s5_ack_i),
    .O(_0193_)
  );
OBUF  _2261_ (
    .I(_0194_[0]),
    .O(s5_addr_o[0])
  );
OBUF  _2262_ (
    .I(_0194_[1]),
    .O(s5_addr_o[1])
  );
OBUF  _2263_ (
    .I(_0194_[10]),
    .O(s5_addr_o[10])
  );
OBUF  _2264_ (
    .I(_0194_[11]),
    .O(s5_addr_o[11])
  );
OBUF  _2265_ (
    .I(_0194_[12]),
    .O(s5_addr_o[12])
  );
OBUF  _2266_ (
    .I(_0194_[13]),
    .O(s5_addr_o[13])
  );
OBUF  _2267_ (
    .I(_0194_[14]),
    .O(s5_addr_o[14])
  );
OBUF  _2268_ (
    .I(_0194_[15]),
    .O(s5_addr_o[15])
  );
OBUF  _2269_ (
    .I(_0194_[16]),
    .O(s5_addr_o[16])
  );
OBUF  _2270_ (
    .I(_0194_[17]),
    .O(s5_addr_o[17])
  );
OBUF  _2271_ (
    .I(_0194_[18]),
    .O(s5_addr_o[18])
  );
OBUF  _2272_ (
    .I(_0194_[19]),
    .O(s5_addr_o[19])
  );
OBUF  _2273_ (
    .I(_0194_[2]),
    .O(s5_addr_o[2])
  );
OBUF  _2274_ (
    .I(_0194_[20]),
    .O(s5_addr_o[20])
  );
OBUF  _2275_ (
    .I(_0194_[21]),
    .O(s5_addr_o[21])
  );
OBUF  _2276_ (
    .I(_0194_[22]),
    .O(s5_addr_o[22])
  );
OBUF  _2277_ (
    .I(_0194_[23]),
    .O(s5_addr_o[23])
  );
OBUF  _2278_ (
    .I(_0194_[24]),
    .O(s5_addr_o[24])
  );
OBUF  _2279_ (
    .I(_0194_[25]),
    .O(s5_addr_o[25])
  );
OBUF  _2280_ (
    .I(_0194_[26]),
    .O(s5_addr_o[26])
  );
OBUF  _2281_ (
    .I(_0194_[27]),
    .O(s5_addr_o[27])
  );
OBUF  _2282_ (
    .I(_0194_[28]),
    .O(s5_addr_o[28])
  );
OBUF  _2283_ (
    .I(_0194_[29]),
    .O(s5_addr_o[29])
  );
OBUF  _2284_ (
    .I(_0194_[3]),
    .O(s5_addr_o[3])
  );
OBUF  _2285_ (
    .I(_0194_[30]),
    .O(s5_addr_o[30])
  );
OBUF  _2286_ (
    .I(_0194_[31]),
    .O(s5_addr_o[31])
  );
OBUF  _2287_ (
    .I(_0194_[4]),
    .O(s5_addr_o[4])
  );
OBUF  _2288_ (
    .I(_0194_[5]),
    .O(s5_addr_o[5])
  );
OBUF  _2289_ (
    .I(_0194_[6]),
    .O(s5_addr_o[6])
  );
OBUF  _2290_ (
    .I(_0194_[7]),
    .O(s5_addr_o[7])
  );
OBUF  _2291_ (
    .I(_0194_[8]),
    .O(s5_addr_o[8])
  );
OBUF  _2292_ (
    .I(_0194_[9]),
    .O(s5_addr_o[9])
  );
OBUF  _2293_ (
    .I(_0195_),
    .O(s5_cyc_o)
  );
IBUF  _2294_ (
    .I(s5_data_i[0]),
    .O(_0196_[0])
  );
IBUF  _2295_ (
    .I(s5_data_i[1]),
    .O(_0196_[1])
  );
IBUF  _2296_ (
    .I(s5_data_i[10]),
    .O(_0196_[10])
  );
IBUF  _2297_ (
    .I(s5_data_i[11]),
    .O(_0196_[11])
  );
IBUF  _2298_ (
    .I(s5_data_i[12]),
    .O(_0196_[12])
  );
IBUF  _2299_ (
    .I(s5_data_i[13]),
    .O(_0196_[13])
  );
IBUF  _2300_ (
    .I(s5_data_i[14]),
    .O(_0196_[14])
  );
IBUF  _2301_ (
    .I(s5_data_i[15]),
    .O(_0196_[15])
  );
IBUF  _2302_ (
    .I(s5_data_i[16]),
    .O(_0196_[16])
  );
IBUF  _2303_ (
    .I(s5_data_i[17]),
    .O(_0196_[17])
  );
IBUF  _2304_ (
    .I(s5_data_i[18]),
    .O(_0196_[18])
  );
IBUF  _2305_ (
    .I(s5_data_i[19]),
    .O(_0196_[19])
  );
IBUF  _2306_ (
    .I(s5_data_i[2]),
    .O(_0196_[2])
  );
IBUF  _2307_ (
    .I(s5_data_i[20]),
    .O(_0196_[20])
  );
IBUF  _2308_ (
    .I(s5_data_i[21]),
    .O(_0196_[21])
  );
IBUF  _2309_ (
    .I(s5_data_i[22]),
    .O(_0196_[22])
  );
IBUF  _2310_ (
    .I(s5_data_i[23]),
    .O(_0196_[23])
  );
IBUF  _2311_ (
    .I(s5_data_i[24]),
    .O(_0196_[24])
  );
IBUF  _2312_ (
    .I(s5_data_i[25]),
    .O(_0196_[25])
  );
IBUF  _2313_ (
    .I(s5_data_i[26]),
    .O(_0196_[26])
  );
IBUF  _2314_ (
    .I(s5_data_i[27]),
    .O(_0196_[27])
  );
IBUF  _2315_ (
    .I(s5_data_i[28]),
    .O(_0196_[28])
  );
IBUF  _2316_ (
    .I(s5_data_i[29]),
    .O(_0196_[29])
  );
IBUF  _2317_ (
    .I(s5_data_i[3]),
    .O(_0196_[3])
  );
IBUF  _2318_ (
    .I(s5_data_i[30]),
    .O(_0196_[30])
  );
IBUF  _2319_ (
    .I(s5_data_i[31]),
    .O(_0196_[31])
  );
IBUF  _2320_ (
    .I(s5_data_i[4]),
    .O(_0196_[4])
  );
IBUF  _2321_ (
    .I(s5_data_i[5]),
    .O(_0196_[5])
  );
IBUF  _2322_ (
    .I(s5_data_i[6]),
    .O(_0196_[6])
  );
IBUF  _2323_ (
    .I(s5_data_i[7]),
    .O(_0196_[7])
  );
IBUF  _2324_ (
    .I(s5_data_i[8]),
    .O(_0196_[8])
  );
IBUF  _2325_ (
    .I(s5_data_i[9]),
    .O(_0196_[9])
  );
OBUF  _2326_ (
    .I(_0197_[0]),
    .O(s5_data_o[0])
  );
OBUF  _2327_ (
    .I(_0197_[1]),
    .O(s5_data_o[1])
  );
OBUF  _2328_ (
    .I(_0197_[10]),
    .O(s5_data_o[10])
  );
OBUF  _2329_ (
    .I(_0197_[11]),
    .O(s5_data_o[11])
  );
OBUF  _2330_ (
    .I(_0197_[12]),
    .O(s5_data_o[12])
  );
OBUF  _2331_ (
    .I(_0197_[13]),
    .O(s5_data_o[13])
  );
OBUF  _2332_ (
    .I(_0197_[14]),
    .O(s5_data_o[14])
  );
OBUF  _2333_ (
    .I(_0197_[15]),
    .O(s5_data_o[15])
  );
OBUF  _2334_ (
    .I(_0197_[16]),
    .O(s5_data_o[16])
  );
OBUF  _2335_ (
    .I(_0197_[17]),
    .O(s5_data_o[17])
  );
OBUF  _2336_ (
    .I(_0197_[18]),
    .O(s5_data_o[18])
  );
OBUF  _2337_ (
    .I(_0197_[19]),
    .O(s5_data_o[19])
  );
OBUF  _2338_ (
    .I(_0197_[2]),
    .O(s5_data_o[2])
  );
OBUF  _2339_ (
    .I(_0197_[20]),
    .O(s5_data_o[20])
  );
OBUF  _2340_ (
    .I(_0197_[21]),
    .O(s5_data_o[21])
  );
OBUF  _2341_ (
    .I(_0197_[22]),
    .O(s5_data_o[22])
  );
OBUF  _2342_ (
    .I(_0197_[23]),
    .O(s5_data_o[23])
  );
OBUF  _2343_ (
    .I(_0197_[24]),
    .O(s5_data_o[24])
  );
OBUF  _2344_ (
    .I(_0197_[25]),
    .O(s5_data_o[25])
  );
OBUF  _2345_ (
    .I(_0197_[26]),
    .O(s5_data_o[26])
  );
OBUF  _2346_ (
    .I(_0197_[27]),
    .O(s5_data_o[27])
  );
OBUF  _2347_ (
    .I(_0197_[28]),
    .O(s5_data_o[28])
  );
OBUF  _2348_ (
    .I(_0197_[29]),
    .O(s5_data_o[29])
  );
OBUF  _2349_ (
    .I(_0197_[3]),
    .O(s5_data_o[3])
  );
OBUF  _2350_ (
    .I(_0197_[30]),
    .O(s5_data_o[30])
  );
OBUF  _2351_ (
    .I(_0197_[31]),
    .O(s5_data_o[31])
  );
OBUF  _2352_ (
    .I(_0197_[4]),
    .O(s5_data_o[4])
  );
OBUF  _2353_ (
    .I(_0197_[5]),
    .O(s5_data_o[5])
  );
OBUF  _2354_ (
    .I(_0197_[6]),
    .O(s5_data_o[6])
  );
OBUF  _2355_ (
    .I(_0197_[7]),
    .O(s5_data_o[7])
  );
OBUF  _2356_ (
    .I(_0197_[8]),
    .O(s5_data_o[8])
  );
OBUF  _2357_ (
    .I(_0197_[9]),
    .O(s5_data_o[9])
  );
IBUF  _2358_ (
    .I(s5_err_i),
    .O(_0198_)
  );
IBUF  _2359_ (
    .I(s5_rty_i),
    .O(_0199_)
  );
OBUF  _2360_ (
    .I(_0200_[0]),
    .O(s5_sel_o[0])
  );
OBUF  _2361_ (
    .I(_0200_[1]),
    .O(s5_sel_o[1])
  );
OBUF  _2362_ (
    .I(_0200_[2]),
    .O(s5_sel_o[2])
  );
OBUF  _2363_ (
    .I(_0200_[3]),
    .O(s5_sel_o[3])
  );
OBUF  _2364_ (
    .I(_0201_),
    .O(s5_stb_o)
  );
OBUF  _2365_ (
    .I(_0202_),
    .O(s5_we_o)
  );
IBUF  _2366_ (
    .I(s6_ack_i),
    .O(_0203_)
  );
OBUF  _2367_ (
    .I(_0204_[0]),
    .O(s6_addr_o[0])
  );
OBUF  _2368_ (
    .I(_0204_[1]),
    .O(s6_addr_o[1])
  );
OBUF  _2369_ (
    .I(_0204_[10]),
    .O(s6_addr_o[10])
  );
OBUF  _2370_ (
    .I(_0204_[11]),
    .O(s6_addr_o[11])
  );
OBUF  _2371_ (
    .I(_0204_[12]),
    .O(s6_addr_o[12])
  );
OBUF  _2372_ (
    .I(_0204_[13]),
    .O(s6_addr_o[13])
  );
OBUF  _2373_ (
    .I(_0204_[14]),
    .O(s6_addr_o[14])
  );
OBUF  _2374_ (
    .I(_0204_[15]),
    .O(s6_addr_o[15])
  );
OBUF  _2375_ (
    .I(_0204_[16]),
    .O(s6_addr_o[16])
  );
OBUF  _2376_ (
    .I(_0204_[17]),
    .O(s6_addr_o[17])
  );
OBUF  _2377_ (
    .I(_0204_[18]),
    .O(s6_addr_o[18])
  );
OBUF  _2378_ (
    .I(_0204_[19]),
    .O(s6_addr_o[19])
  );
OBUF  _2379_ (
    .I(_0204_[2]),
    .O(s6_addr_o[2])
  );
OBUF  _2380_ (
    .I(_0204_[20]),
    .O(s6_addr_o[20])
  );
OBUF  _2381_ (
    .I(_0204_[21]),
    .O(s6_addr_o[21])
  );
OBUF  _2382_ (
    .I(_0204_[22]),
    .O(s6_addr_o[22])
  );
OBUF  _2383_ (
    .I(_0204_[23]),
    .O(s6_addr_o[23])
  );
OBUF  _2384_ (
    .I(_0204_[24]),
    .O(s6_addr_o[24])
  );
OBUF  _2385_ (
    .I(_0204_[25]),
    .O(s6_addr_o[25])
  );
OBUF  _2386_ (
    .I(_0204_[26]),
    .O(s6_addr_o[26])
  );
OBUF  _2387_ (
    .I(_0204_[27]),
    .O(s6_addr_o[27])
  );
OBUF  _2388_ (
    .I(_0204_[28]),
    .O(s6_addr_o[28])
  );
OBUF  _2389_ (
    .I(_0204_[29]),
    .O(s6_addr_o[29])
  );
OBUF  _2390_ (
    .I(_0204_[3]),
    .O(s6_addr_o[3])
  );
OBUF  _2391_ (
    .I(_0204_[30]),
    .O(s6_addr_o[30])
  );
OBUF  _2392_ (
    .I(_0204_[31]),
    .O(s6_addr_o[31])
  );
OBUF  _2393_ (
    .I(_0204_[4]),
    .O(s6_addr_o[4])
  );
OBUF  _2394_ (
    .I(_0204_[5]),
    .O(s6_addr_o[5])
  );
OBUF  _2395_ (
    .I(_0204_[6]),
    .O(s6_addr_o[6])
  );
OBUF  _2396_ (
    .I(_0204_[7]),
    .O(s6_addr_o[7])
  );
OBUF  _2397_ (
    .I(_0204_[8]),
    .O(s6_addr_o[8])
  );
OBUF  _2398_ (
    .I(_0204_[9]),
    .O(s6_addr_o[9])
  );
OBUF  _2399_ (
    .I(_0205_),
    .O(s6_cyc_o)
  );
IBUF  _2400_ (
    .I(s6_data_i[0]),
    .O(_0206_[0])
  );
IBUF  _2401_ (
    .I(s6_data_i[1]),
    .O(_0206_[1])
  );
IBUF  _2402_ (
    .I(s6_data_i[10]),
    .O(_0206_[10])
  );
IBUF  _2403_ (
    .I(s6_data_i[11]),
    .O(_0206_[11])
  );
IBUF  _2404_ (
    .I(s6_data_i[12]),
    .O(_0206_[12])
  );
IBUF  _2405_ (
    .I(s6_data_i[13]),
    .O(_0206_[13])
  );
IBUF  _2406_ (
    .I(s6_data_i[14]),
    .O(_0206_[14])
  );
IBUF  _2407_ (
    .I(s6_data_i[15]),
    .O(_0206_[15])
  );
IBUF  _2408_ (
    .I(s6_data_i[16]),
    .O(_0206_[16])
  );
IBUF  _2409_ (
    .I(s6_data_i[17]),
    .O(_0206_[17])
  );
IBUF  _2410_ (
    .I(s6_data_i[18]),
    .O(_0206_[18])
  );
IBUF  _2411_ (
    .I(s6_data_i[19]),
    .O(_0206_[19])
  );
IBUF  _2412_ (
    .I(s6_data_i[2]),
    .O(_0206_[2])
  );
IBUF  _2413_ (
    .I(s6_data_i[20]),
    .O(_0206_[20])
  );
IBUF  _2414_ (
    .I(s6_data_i[21]),
    .O(_0206_[21])
  );
IBUF  _2415_ (
    .I(s6_data_i[22]),
    .O(_0206_[22])
  );
IBUF  _2416_ (
    .I(s6_data_i[23]),
    .O(_0206_[23])
  );
IBUF  _2417_ (
    .I(s6_data_i[24]),
    .O(_0206_[24])
  );
IBUF  _2418_ (
    .I(s6_data_i[25]),
    .O(_0206_[25])
  );
IBUF  _2419_ (
    .I(s6_data_i[26]),
    .O(_0206_[26])
  );
IBUF  _2420_ (
    .I(s6_data_i[27]),
    .O(_0206_[27])
  );
IBUF  _2421_ (
    .I(s6_data_i[28]),
    .O(_0206_[28])
  );
IBUF  _2422_ (
    .I(s6_data_i[29]),
    .O(_0206_[29])
  );
IBUF  _2423_ (
    .I(s6_data_i[3]),
    .O(_0206_[3])
  );
IBUF  _2424_ (
    .I(s6_data_i[30]),
    .O(_0206_[30])
  );
IBUF  _2425_ (
    .I(s6_data_i[31]),
    .O(_0206_[31])
  );
IBUF  _2426_ (
    .I(s6_data_i[4]),
    .O(_0206_[4])
  );
IBUF  _2427_ (
    .I(s6_data_i[5]),
    .O(_0206_[5])
  );
IBUF  _2428_ (
    .I(s6_data_i[6]),
    .O(_0206_[6])
  );
IBUF  _2429_ (
    .I(s6_data_i[7]),
    .O(_0206_[7])
  );
IBUF  _2430_ (
    .I(s6_data_i[8]),
    .O(_0206_[8])
  );
IBUF  _2431_ (
    .I(s6_data_i[9]),
    .O(_0206_[9])
  );
OBUF  _2432_ (
    .I(_0207_[0]),
    .O(s6_data_o[0])
  );
OBUF  _2433_ (
    .I(_0207_[1]),
    .O(s6_data_o[1])
  );
OBUF  _2434_ (
    .I(_0207_[10]),
    .O(s6_data_o[10])
  );
OBUF  _2435_ (
    .I(_0207_[11]),
    .O(s6_data_o[11])
  );
OBUF  _2436_ (
    .I(_0207_[12]),
    .O(s6_data_o[12])
  );
OBUF  _2437_ (
    .I(_0207_[13]),
    .O(s6_data_o[13])
  );
OBUF  _2438_ (
    .I(_0207_[14]),
    .O(s6_data_o[14])
  );
OBUF  _2439_ (
    .I(_0207_[15]),
    .O(s6_data_o[15])
  );
OBUF  _2440_ (
    .I(_0207_[16]),
    .O(s6_data_o[16])
  );
OBUF  _2441_ (
    .I(_0207_[17]),
    .O(s6_data_o[17])
  );
OBUF  _2442_ (
    .I(_0207_[18]),
    .O(s6_data_o[18])
  );
OBUF  _2443_ (
    .I(_0207_[19]),
    .O(s6_data_o[19])
  );
OBUF  _2444_ (
    .I(_0207_[2]),
    .O(s6_data_o[2])
  );
OBUF  _2445_ (
    .I(_0207_[20]),
    .O(s6_data_o[20])
  );
OBUF  _2446_ (
    .I(_0207_[21]),
    .O(s6_data_o[21])
  );
OBUF  _2447_ (
    .I(_0207_[22]),
    .O(s6_data_o[22])
  );
OBUF  _2448_ (
    .I(_0207_[23]),
    .O(s6_data_o[23])
  );
OBUF  _2449_ (
    .I(_0207_[24]),
    .O(s6_data_o[24])
  );
OBUF  _2450_ (
    .I(_0207_[25]),
    .O(s6_data_o[25])
  );
OBUF  _2451_ (
    .I(_0207_[26]),
    .O(s6_data_o[26])
  );
OBUF  _2452_ (
    .I(_0207_[27]),
    .O(s6_data_o[27])
  );
OBUF  _2453_ (
    .I(_0207_[28]),
    .O(s6_data_o[28])
  );
OBUF  _2454_ (
    .I(_0207_[29]),
    .O(s6_data_o[29])
  );
OBUF  _2455_ (
    .I(_0207_[3]),
    .O(s6_data_o[3])
  );
OBUF  _2456_ (
    .I(_0207_[30]),
    .O(s6_data_o[30])
  );
OBUF  _2457_ (
    .I(_0207_[31]),
    .O(s6_data_o[31])
  );
OBUF  _2458_ (
    .I(_0207_[4]),
    .O(s6_data_o[4])
  );
OBUF  _2459_ (
    .I(_0207_[5]),
    .O(s6_data_o[5])
  );
OBUF  _2460_ (
    .I(_0207_[6]),
    .O(s6_data_o[6])
  );
OBUF  _2461_ (
    .I(_0207_[7]),
    .O(s6_data_o[7])
  );
OBUF  _2462_ (
    .I(_0207_[8]),
    .O(s6_data_o[8])
  );
OBUF  _2463_ (
    .I(_0207_[9]),
    .O(s6_data_o[9])
  );
IBUF  _2464_ (
    .I(s6_err_i),
    .O(_0208_)
  );
IBUF  _2465_ (
    .I(s6_rty_i),
    .O(_0209_)
  );
OBUF  _2466_ (
    .I(_0210_[0]),
    .O(s6_sel_o[0])
  );
OBUF  _2467_ (
    .I(_0210_[1]),
    .O(s6_sel_o[1])
  );
OBUF  _2468_ (
    .I(_0210_[2]),
    .O(s6_sel_o[2])
  );
OBUF  _2469_ (
    .I(_0210_[3]),
    .O(s6_sel_o[3])
  );
OBUF  _2470_ (
    .I(_0211_),
    .O(s6_stb_o)
  );
OBUF  _2471_ (
    .I(_0212_),
    .O(s6_we_o)
  );
IBUF  _2472_ (
    .I(s7_ack_i),
    .O(_0213_)
  );
OBUF  _2473_ (
    .I(_0214_[0]),
    .O(s7_addr_o[0])
  );
OBUF  _2474_ (
    .I(_0214_[1]),
    .O(s7_addr_o[1])
  );
OBUF  _2475_ (
    .I(_0214_[10]),
    .O(s7_addr_o[10])
  );
OBUF  _2476_ (
    .I(_0214_[11]),
    .O(s7_addr_o[11])
  );
OBUF  _2477_ (
    .I(_0214_[12]),
    .O(s7_addr_o[12])
  );
OBUF  _2478_ (
    .I(_0214_[13]),
    .O(s7_addr_o[13])
  );
OBUF  _2479_ (
    .I(_0214_[14]),
    .O(s7_addr_o[14])
  );
OBUF  _2480_ (
    .I(_0214_[15]),
    .O(s7_addr_o[15])
  );
OBUF  _2481_ (
    .I(_0214_[16]),
    .O(s7_addr_o[16])
  );
OBUF  _2482_ (
    .I(_0214_[17]),
    .O(s7_addr_o[17])
  );
OBUF  _2483_ (
    .I(_0214_[18]),
    .O(s7_addr_o[18])
  );
OBUF  _2484_ (
    .I(_0214_[19]),
    .O(s7_addr_o[19])
  );
OBUF  _2485_ (
    .I(_0214_[2]),
    .O(s7_addr_o[2])
  );
OBUF  _2486_ (
    .I(_0214_[20]),
    .O(s7_addr_o[20])
  );
OBUF  _2487_ (
    .I(_0214_[21]),
    .O(s7_addr_o[21])
  );
OBUF  _2488_ (
    .I(_0214_[22]),
    .O(s7_addr_o[22])
  );
OBUF  _2489_ (
    .I(_0214_[23]),
    .O(s7_addr_o[23])
  );
OBUF  _2490_ (
    .I(_0214_[24]),
    .O(s7_addr_o[24])
  );
OBUF  _2491_ (
    .I(_0214_[25]),
    .O(s7_addr_o[25])
  );
OBUF  _2492_ (
    .I(_0214_[26]),
    .O(s7_addr_o[26])
  );
OBUF  _2493_ (
    .I(_0214_[27]),
    .O(s7_addr_o[27])
  );
OBUF  _2494_ (
    .I(_0214_[28]),
    .O(s7_addr_o[28])
  );
OBUF  _2495_ (
    .I(_0214_[29]),
    .O(s7_addr_o[29])
  );
OBUF  _2496_ (
    .I(_0214_[3]),
    .O(s7_addr_o[3])
  );
OBUF  _2497_ (
    .I(_0214_[30]),
    .O(s7_addr_o[30])
  );
OBUF  _2498_ (
    .I(_0214_[31]),
    .O(s7_addr_o[31])
  );
OBUF  _2499_ (
    .I(_0214_[4]),
    .O(s7_addr_o[4])
  );
OBUF  _2500_ (
    .I(_0214_[5]),
    .O(s7_addr_o[5])
  );
OBUF  _2501_ (
    .I(_0214_[6]),
    .O(s7_addr_o[6])
  );
OBUF  _2502_ (
    .I(_0214_[7]),
    .O(s7_addr_o[7])
  );
OBUF  _2503_ (
    .I(_0214_[8]),
    .O(s7_addr_o[8])
  );
OBUF  _2504_ (
    .I(_0214_[9]),
    .O(s7_addr_o[9])
  );
OBUF  _2505_ (
    .I(_0215_),
    .O(s7_cyc_o)
  );
IBUF  _2506_ (
    .I(s7_data_i[0]),
    .O(_0216_[0])
  );
IBUF  _2507_ (
    .I(s7_data_i[1]),
    .O(_0216_[1])
  );
IBUF  _2508_ (
    .I(s7_data_i[10]),
    .O(_0216_[10])
  );
IBUF  _2509_ (
    .I(s7_data_i[11]),
    .O(_0216_[11])
  );
IBUF  _2510_ (
    .I(s7_data_i[12]),
    .O(_0216_[12])
  );
IBUF  _2511_ (
    .I(s7_data_i[13]),
    .O(_0216_[13])
  );
IBUF  _2512_ (
    .I(s7_data_i[14]),
    .O(_0216_[14])
  );
IBUF  _2513_ (
    .I(s7_data_i[15]),
    .O(_0216_[15])
  );
IBUF  _2514_ (
    .I(s7_data_i[16]),
    .O(_0216_[16])
  );
IBUF  _2515_ (
    .I(s7_data_i[17]),
    .O(_0216_[17])
  );
IBUF  _2516_ (
    .I(s7_data_i[18]),
    .O(_0216_[18])
  );
IBUF  _2517_ (
    .I(s7_data_i[19]),
    .O(_0216_[19])
  );
IBUF  _2518_ (
    .I(s7_data_i[2]),
    .O(_0216_[2])
  );
IBUF  _2519_ (
    .I(s7_data_i[20]),
    .O(_0216_[20])
  );
IBUF  _2520_ (
    .I(s7_data_i[21]),
    .O(_0216_[21])
  );
IBUF  _2521_ (
    .I(s7_data_i[22]),
    .O(_0216_[22])
  );
IBUF  _2522_ (
    .I(s7_data_i[23]),
    .O(_0216_[23])
  );
IBUF  _2523_ (
    .I(s7_data_i[24]),
    .O(_0216_[24])
  );
IBUF  _2524_ (
    .I(s7_data_i[25]),
    .O(_0216_[25])
  );
IBUF  _2525_ (
    .I(s7_data_i[26]),
    .O(_0216_[26])
  );
IBUF  _2526_ (
    .I(s7_data_i[27]),
    .O(_0216_[27])
  );
IBUF  _2527_ (
    .I(s7_data_i[28]),
    .O(_0216_[28])
  );
IBUF  _2528_ (
    .I(s7_data_i[29]),
    .O(_0216_[29])
  );
IBUF  _2529_ (
    .I(s7_data_i[3]),
    .O(_0216_[3])
  );
IBUF  _2530_ (
    .I(s7_data_i[30]),
    .O(_0216_[30])
  );
IBUF  _2531_ (
    .I(s7_data_i[31]),
    .O(_0216_[31])
  );
IBUF  _2532_ (
    .I(s7_data_i[4]),
    .O(_0216_[4])
  );
IBUF  _2533_ (
    .I(s7_data_i[5]),
    .O(_0216_[5])
  );
IBUF  _2534_ (
    .I(s7_data_i[6]),
    .O(_0216_[6])
  );
IBUF  _2535_ (
    .I(s7_data_i[7]),
    .O(_0216_[7])
  );
IBUF  _2536_ (
    .I(s7_data_i[8]),
    .O(_0216_[8])
  );
IBUF  _2537_ (
    .I(s7_data_i[9]),
    .O(_0216_[9])
  );
OBUF  _2538_ (
    .I(_0217_[0]),
    .O(s7_data_o[0])
  );
OBUF  _2539_ (
    .I(_0217_[1]),
    .O(s7_data_o[1])
  );
OBUF  _2540_ (
    .I(_0217_[10]),
    .O(s7_data_o[10])
  );
OBUF  _2541_ (
    .I(_0217_[11]),
    .O(s7_data_o[11])
  );
OBUF  _2542_ (
    .I(_0217_[12]),
    .O(s7_data_o[12])
  );
OBUF  _2543_ (
    .I(_0217_[13]),
    .O(s7_data_o[13])
  );
OBUF  _2544_ (
    .I(_0217_[14]),
    .O(s7_data_o[14])
  );
OBUF  _2545_ (
    .I(_0217_[15]),
    .O(s7_data_o[15])
  );
OBUF  _2546_ (
    .I(_0217_[16]),
    .O(s7_data_o[16])
  );
OBUF  _2547_ (
    .I(_0217_[17]),
    .O(s7_data_o[17])
  );
OBUF  _2548_ (
    .I(_0217_[18]),
    .O(s7_data_o[18])
  );
OBUF  _2549_ (
    .I(_0217_[19]),
    .O(s7_data_o[19])
  );
OBUF  _2550_ (
    .I(_0217_[2]),
    .O(s7_data_o[2])
  );
OBUF  _2551_ (
    .I(_0217_[20]),
    .O(s7_data_o[20])
  );
OBUF  _2552_ (
    .I(_0217_[21]),
    .O(s7_data_o[21])
  );
OBUF  _2553_ (
    .I(_0217_[22]),
    .O(s7_data_o[22])
  );
OBUF  _2554_ (
    .I(_0217_[23]),
    .O(s7_data_o[23])
  );
OBUF  _2555_ (
    .I(_0217_[24]),
    .O(s7_data_o[24])
  );
OBUF  _2556_ (
    .I(_0217_[25]),
    .O(s7_data_o[25])
  );
OBUF  _2557_ (
    .I(_0217_[26]),
    .O(s7_data_o[26])
  );
OBUF  _2558_ (
    .I(_0217_[27]),
    .O(s7_data_o[27])
  );
OBUF  _2559_ (
    .I(_0217_[28]),
    .O(s7_data_o[28])
  );
OBUF  _2560_ (
    .I(_0217_[29]),
    .O(s7_data_o[29])
  );
OBUF  _2561_ (
    .I(_0217_[3]),
    .O(s7_data_o[3])
  );
OBUF  _2562_ (
    .I(_0217_[30]),
    .O(s7_data_o[30])
  );
OBUF  _2563_ (
    .I(_0217_[31]),
    .O(s7_data_o[31])
  );
OBUF  _2564_ (
    .I(_0217_[4]),
    .O(s7_data_o[4])
  );
OBUF  _2565_ (
    .I(_0217_[5]),
    .O(s7_data_o[5])
  );
OBUF  _2566_ (
    .I(_0217_[6]),
    .O(s7_data_o[6])
  );
OBUF  _2567_ (
    .I(_0217_[7]),
    .O(s7_data_o[7])
  );
OBUF  _2568_ (
    .I(_0217_[8]),
    .O(s7_data_o[8])
  );
OBUF  _2569_ (
    .I(_0217_[9]),
    .O(s7_data_o[9])
  );
IBUF  _2570_ (
    .I(s7_err_i),
    .O(_0218_)
  );
IBUF  _2571_ (
    .I(s7_rty_i),
    .O(_0219_)
  );
OBUF  _2572_ (
    .I(_0220_[0]),
    .O(s7_sel_o[0])
  );
OBUF  _2573_ (
    .I(_0220_[1]),
    .O(s7_sel_o[1])
  );
OBUF  _2574_ (
    .I(_0220_[2]),
    .O(s7_sel_o[2])
  );
OBUF  _2575_ (
    .I(_0220_[3]),
    .O(s7_sel_o[3])
  );
OBUF  _2576_ (
    .I(_0221_),
    .O(s7_stb_o)
  );
OBUF  _2577_ (
    .I(_0222_),
    .O(s7_we_o)
  );
IBUF  _2578_ (
    .I(s8_ack_i),
    .O(_0223_)
  );
OBUF  _2579_ (
    .I(_0224_[0]),
    .O(s8_addr_o[0])
  );
OBUF  _2580_ (
    .I(_0224_[1]),
    .O(s8_addr_o[1])
  );
OBUF  _2581_ (
    .I(_0224_[10]),
    .O(s8_addr_o[10])
  );
OBUF  _2582_ (
    .I(_0224_[11]),
    .O(s8_addr_o[11])
  );
OBUF  _2583_ (
    .I(_0224_[12]),
    .O(s8_addr_o[12])
  );
OBUF  _2584_ (
    .I(_0224_[13]),
    .O(s8_addr_o[13])
  );
OBUF  _2585_ (
    .I(_0224_[14]),
    .O(s8_addr_o[14])
  );
OBUF  _2586_ (
    .I(_0224_[15]),
    .O(s8_addr_o[15])
  );
OBUF  _2587_ (
    .I(_0224_[16]),
    .O(s8_addr_o[16])
  );
OBUF  _2588_ (
    .I(_0224_[17]),
    .O(s8_addr_o[17])
  );
OBUF  _2589_ (
    .I(_0224_[18]),
    .O(s8_addr_o[18])
  );
OBUF  _2590_ (
    .I(_0224_[19]),
    .O(s8_addr_o[19])
  );
OBUF  _2591_ (
    .I(_0224_[2]),
    .O(s8_addr_o[2])
  );
OBUF  _2592_ (
    .I(_0224_[20]),
    .O(s8_addr_o[20])
  );
OBUF  _2593_ (
    .I(_0224_[21]),
    .O(s8_addr_o[21])
  );
OBUF  _2594_ (
    .I(_0224_[22]),
    .O(s8_addr_o[22])
  );
OBUF  _2595_ (
    .I(_0224_[23]),
    .O(s8_addr_o[23])
  );
OBUF  _2596_ (
    .I(_0224_[24]),
    .O(s8_addr_o[24])
  );
OBUF  _2597_ (
    .I(_0224_[25]),
    .O(s8_addr_o[25])
  );
OBUF  _2598_ (
    .I(_0224_[26]),
    .O(s8_addr_o[26])
  );
OBUF  _2599_ (
    .I(_0224_[27]),
    .O(s8_addr_o[27])
  );
OBUF  _2600_ (
    .I(_0224_[28]),
    .O(s8_addr_o[28])
  );
OBUF  _2601_ (
    .I(_0224_[29]),
    .O(s8_addr_o[29])
  );
OBUF  _2602_ (
    .I(_0224_[3]),
    .O(s8_addr_o[3])
  );
OBUF  _2603_ (
    .I(_0224_[30]),
    .O(s8_addr_o[30])
  );
OBUF  _2604_ (
    .I(_0224_[31]),
    .O(s8_addr_o[31])
  );
OBUF  _2605_ (
    .I(_0224_[4]),
    .O(s8_addr_o[4])
  );
OBUF  _2606_ (
    .I(_0224_[5]),
    .O(s8_addr_o[5])
  );
OBUF  _2607_ (
    .I(_0224_[6]),
    .O(s8_addr_o[6])
  );
OBUF  _2608_ (
    .I(_0224_[7]),
    .O(s8_addr_o[7])
  );
OBUF  _2609_ (
    .I(_0224_[8]),
    .O(s8_addr_o[8])
  );
OBUF  _2610_ (
    .I(_0224_[9]),
    .O(s8_addr_o[9])
  );
OBUF  _2611_ (
    .I(_0225_),
    .O(s8_cyc_o)
  );
IBUF  _2612_ (
    .I(s8_data_i[0]),
    .O(_0226_[0])
  );
IBUF  _2613_ (
    .I(s8_data_i[1]),
    .O(_0226_[1])
  );
IBUF  _2614_ (
    .I(s8_data_i[10]),
    .O(_0226_[10])
  );
IBUF  _2615_ (
    .I(s8_data_i[11]),
    .O(_0226_[11])
  );
IBUF  _2616_ (
    .I(s8_data_i[12]),
    .O(_0226_[12])
  );
IBUF  _2617_ (
    .I(s8_data_i[13]),
    .O(_0226_[13])
  );
IBUF  _2618_ (
    .I(s8_data_i[14]),
    .O(_0226_[14])
  );
IBUF  _2619_ (
    .I(s8_data_i[15]),
    .O(_0226_[15])
  );
IBUF  _2620_ (
    .I(s8_data_i[16]),
    .O(_0226_[16])
  );
IBUF  _2621_ (
    .I(s8_data_i[17]),
    .O(_0226_[17])
  );
IBUF  _2622_ (
    .I(s8_data_i[18]),
    .O(_0226_[18])
  );
IBUF  _2623_ (
    .I(s8_data_i[19]),
    .O(_0226_[19])
  );
IBUF  _2624_ (
    .I(s8_data_i[2]),
    .O(_0226_[2])
  );
IBUF  _2625_ (
    .I(s8_data_i[20]),
    .O(_0226_[20])
  );
IBUF  _2626_ (
    .I(s8_data_i[21]),
    .O(_0226_[21])
  );
IBUF  _2627_ (
    .I(s8_data_i[22]),
    .O(_0226_[22])
  );
IBUF  _2628_ (
    .I(s8_data_i[23]),
    .O(_0226_[23])
  );
IBUF  _2629_ (
    .I(s8_data_i[24]),
    .O(_0226_[24])
  );
IBUF  _2630_ (
    .I(s8_data_i[25]),
    .O(_0226_[25])
  );
IBUF  _2631_ (
    .I(s8_data_i[26]),
    .O(_0226_[26])
  );
IBUF  _2632_ (
    .I(s8_data_i[27]),
    .O(_0226_[27])
  );
IBUF  _2633_ (
    .I(s8_data_i[28]),
    .O(_0226_[28])
  );
IBUF  _2634_ (
    .I(s8_data_i[29]),
    .O(_0226_[29])
  );
IBUF  _2635_ (
    .I(s8_data_i[3]),
    .O(_0226_[3])
  );
IBUF  _2636_ (
    .I(s8_data_i[30]),
    .O(_0226_[30])
  );
IBUF  _2637_ (
    .I(s8_data_i[31]),
    .O(_0226_[31])
  );
IBUF  _2638_ (
    .I(s8_data_i[4]),
    .O(_0226_[4])
  );
IBUF  _2639_ (
    .I(s8_data_i[5]),
    .O(_0226_[5])
  );
IBUF  _2640_ (
    .I(s8_data_i[6]),
    .O(_0226_[6])
  );
IBUF  _2641_ (
    .I(s8_data_i[7]),
    .O(_0226_[7])
  );
IBUF  _2642_ (
    .I(s8_data_i[8]),
    .O(_0226_[8])
  );
IBUF  _2643_ (
    .I(s8_data_i[9]),
    .O(_0226_[9])
  );
OBUF  _2644_ (
    .I(_0227_[0]),
    .O(s8_data_o[0])
  );
OBUF  _2645_ (
    .I(_0227_[1]),
    .O(s8_data_o[1])
  );
OBUF  _2646_ (
    .I(_0227_[10]),
    .O(s8_data_o[10])
  );
OBUF  _2647_ (
    .I(_0227_[11]),
    .O(s8_data_o[11])
  );
OBUF  _2648_ (
    .I(_0227_[12]),
    .O(s8_data_o[12])
  );
OBUF  _2649_ (
    .I(_0227_[13]),
    .O(s8_data_o[13])
  );
OBUF  _2650_ (
    .I(_0227_[14]),
    .O(s8_data_o[14])
  );
OBUF  _2651_ (
    .I(_0227_[15]),
    .O(s8_data_o[15])
  );
OBUF  _2652_ (
    .I(_0227_[16]),
    .O(s8_data_o[16])
  );
OBUF  _2653_ (
    .I(_0227_[17]),
    .O(s8_data_o[17])
  );
OBUF  _2654_ (
    .I(_0227_[18]),
    .O(s8_data_o[18])
  );
OBUF  _2655_ (
    .I(_0227_[19]),
    .O(s8_data_o[19])
  );
OBUF  _2656_ (
    .I(_0227_[2]),
    .O(s8_data_o[2])
  );
OBUF  _2657_ (
    .I(_0227_[20]),
    .O(s8_data_o[20])
  );
OBUF  _2658_ (
    .I(_0227_[21]),
    .O(s8_data_o[21])
  );
OBUF  _2659_ (
    .I(_0227_[22]),
    .O(s8_data_o[22])
  );
OBUF  _2660_ (
    .I(_0227_[23]),
    .O(s8_data_o[23])
  );
OBUF  _2661_ (
    .I(_0227_[24]),
    .O(s8_data_o[24])
  );
OBUF  _2662_ (
    .I(_0227_[25]),
    .O(s8_data_o[25])
  );
OBUF  _2663_ (
    .I(_0227_[26]),
    .O(s8_data_o[26])
  );
OBUF  _2664_ (
    .I(_0227_[27]),
    .O(s8_data_o[27])
  );
OBUF  _2665_ (
    .I(_0227_[28]),
    .O(s8_data_o[28])
  );
OBUF  _2666_ (
    .I(_0227_[29]),
    .O(s8_data_o[29])
  );
OBUF  _2667_ (
    .I(_0227_[3]),
    .O(s8_data_o[3])
  );
OBUF  _2668_ (
    .I(_0227_[30]),
    .O(s8_data_o[30])
  );
OBUF  _2669_ (
    .I(_0227_[31]),
    .O(s8_data_o[31])
  );
OBUF  _2670_ (
    .I(_0227_[4]),
    .O(s8_data_o[4])
  );
OBUF  _2671_ (
    .I(_0227_[5]),
    .O(s8_data_o[5])
  );
OBUF  _2672_ (
    .I(_0227_[6]),
    .O(s8_data_o[6])
  );
OBUF  _2673_ (
    .I(_0227_[7]),
    .O(s8_data_o[7])
  );
OBUF  _2674_ (
    .I(_0227_[8]),
    .O(s8_data_o[8])
  );
OBUF  _2675_ (
    .I(_0227_[9]),
    .O(s8_data_o[9])
  );
IBUF  _2676_ (
    .I(s8_err_i),
    .O(_0228_)
  );
IBUF  _2677_ (
    .I(s8_rty_i),
    .O(_0229_)
  );
OBUF  _2678_ (
    .I(_0230_[0]),
    .O(s8_sel_o[0])
  );
OBUF  _2679_ (
    .I(_0230_[1]),
    .O(s8_sel_o[1])
  );
OBUF  _2680_ (
    .I(_0230_[2]),
    .O(s8_sel_o[2])
  );
OBUF  _2681_ (
    .I(_0230_[3]),
    .O(s8_sel_o[3])
  );
OBUF  _2682_ (
    .I(_0231_),
    .O(s8_stb_o)
  );
OBUF  _2683_ (
    .I(_0232_),
    .O(s8_we_o)
  );
IBUF  _2684_ (
    .I(s9_ack_i),
    .O(_0233_)
  );
OBUF  _2685_ (
    .I(_0234_[0]),
    .O(s9_addr_o[0])
  );
OBUF  _2686_ (
    .I(_0234_[1]),
    .O(s9_addr_o[1])
  );
OBUF  _2687_ (
    .I(_0234_[10]),
    .O(s9_addr_o[10])
  );
OBUF  _2688_ (
    .I(_0234_[11]),
    .O(s9_addr_o[11])
  );
OBUF  _2689_ (
    .I(_0234_[12]),
    .O(s9_addr_o[12])
  );
OBUF  _2690_ (
    .I(_0234_[13]),
    .O(s9_addr_o[13])
  );
OBUF  _2691_ (
    .I(_0234_[14]),
    .O(s9_addr_o[14])
  );
OBUF  _2692_ (
    .I(_0234_[15]),
    .O(s9_addr_o[15])
  );
OBUF  _2693_ (
    .I(_0234_[16]),
    .O(s9_addr_o[16])
  );
OBUF  _2694_ (
    .I(_0234_[17]),
    .O(s9_addr_o[17])
  );
OBUF  _2695_ (
    .I(_0234_[18]),
    .O(s9_addr_o[18])
  );
OBUF  _2696_ (
    .I(_0234_[19]),
    .O(s9_addr_o[19])
  );
OBUF  _2697_ (
    .I(_0234_[2]),
    .O(s9_addr_o[2])
  );
OBUF  _2698_ (
    .I(_0234_[20]),
    .O(s9_addr_o[20])
  );
OBUF  _2699_ (
    .I(_0234_[21]),
    .O(s9_addr_o[21])
  );
OBUF  _2700_ (
    .I(_0234_[22]),
    .O(s9_addr_o[22])
  );
OBUF  _2701_ (
    .I(_0234_[23]),
    .O(s9_addr_o[23])
  );
OBUF  _2702_ (
    .I(_0234_[24]),
    .O(s9_addr_o[24])
  );
OBUF  _2703_ (
    .I(_0234_[25]),
    .O(s9_addr_o[25])
  );
OBUF  _2704_ (
    .I(_0234_[26]),
    .O(s9_addr_o[26])
  );
OBUF  _2705_ (
    .I(_0234_[27]),
    .O(s9_addr_o[27])
  );
OBUF  _2706_ (
    .I(_0234_[28]),
    .O(s9_addr_o[28])
  );
OBUF  _2707_ (
    .I(_0234_[29]),
    .O(s9_addr_o[29])
  );
OBUF  _2708_ (
    .I(_0234_[3]),
    .O(s9_addr_o[3])
  );
OBUF  _2709_ (
    .I(_0234_[30]),
    .O(s9_addr_o[30])
  );
OBUF  _2710_ (
    .I(_0234_[31]),
    .O(s9_addr_o[31])
  );
OBUF  _2711_ (
    .I(_0234_[4]),
    .O(s9_addr_o[4])
  );
OBUF  _2712_ (
    .I(_0234_[5]),
    .O(s9_addr_o[5])
  );
OBUF  _2713_ (
    .I(_0234_[6]),
    .O(s9_addr_o[6])
  );
OBUF  _2714_ (
    .I(_0234_[7]),
    .O(s9_addr_o[7])
  );
OBUF  _2715_ (
    .I(_0234_[8]),
    .O(s9_addr_o[8])
  );
OBUF  _2716_ (
    .I(_0234_[9]),
    .O(s9_addr_o[9])
  );
OBUF  _2717_ (
    .I(_0235_),
    .O(s9_cyc_o)
  );
IBUF  _2718_ (
    .I(s9_data_i[0]),
    .O(_0236_[0])
  );
IBUF  _2719_ (
    .I(s9_data_i[1]),
    .O(_0236_[1])
  );
IBUF  _2720_ (
    .I(s9_data_i[10]),
    .O(_0236_[10])
  );
IBUF  _2721_ (
    .I(s9_data_i[11]),
    .O(_0236_[11])
  );
IBUF  _2722_ (
    .I(s9_data_i[12]),
    .O(_0236_[12])
  );
IBUF  _2723_ (
    .I(s9_data_i[13]),
    .O(_0236_[13])
  );
IBUF  _2724_ (
    .I(s9_data_i[14]),
    .O(_0236_[14])
  );
IBUF  _2725_ (
    .I(s9_data_i[15]),
    .O(_0236_[15])
  );
IBUF  _2726_ (
    .I(s9_data_i[16]),
    .O(_0236_[16])
  );
IBUF  _2727_ (
    .I(s9_data_i[17]),
    .O(_0236_[17])
  );
IBUF  _2728_ (
    .I(s9_data_i[18]),
    .O(_0236_[18])
  );
IBUF  _2729_ (
    .I(s9_data_i[19]),
    .O(_0236_[19])
  );
IBUF  _2730_ (
    .I(s9_data_i[2]),
    .O(_0236_[2])
  );
IBUF  _2731_ (
    .I(s9_data_i[20]),
    .O(_0236_[20])
  );
IBUF  _2732_ (
    .I(s9_data_i[21]),
    .O(_0236_[21])
  );
IBUF  _2733_ (
    .I(s9_data_i[22]),
    .O(_0236_[22])
  );
IBUF  _2734_ (
    .I(s9_data_i[23]),
    .O(_0236_[23])
  );
IBUF  _2735_ (
    .I(s9_data_i[24]),
    .O(_0236_[24])
  );
IBUF  _2736_ (
    .I(s9_data_i[25]),
    .O(_0236_[25])
  );
IBUF  _2737_ (
    .I(s9_data_i[26]),
    .O(_0236_[26])
  );
IBUF  _2738_ (
    .I(s9_data_i[27]),
    .O(_0236_[27])
  );
IBUF  _2739_ (
    .I(s9_data_i[28]),
    .O(_0236_[28])
  );
IBUF  _2740_ (
    .I(s9_data_i[29]),
    .O(_0236_[29])
  );
IBUF  _2741_ (
    .I(s9_data_i[3]),
    .O(_0236_[3])
  );
IBUF  _2742_ (
    .I(s9_data_i[30]),
    .O(_0236_[30])
  );
IBUF  _2743_ (
    .I(s9_data_i[31]),
    .O(_0236_[31])
  );
IBUF  _2744_ (
    .I(s9_data_i[4]),
    .O(_0236_[4])
  );
IBUF  _2745_ (
    .I(s9_data_i[5]),
    .O(_0236_[5])
  );
IBUF  _2746_ (
    .I(s9_data_i[6]),
    .O(_0236_[6])
  );
IBUF  _2747_ (
    .I(s9_data_i[7]),
    .O(_0236_[7])
  );
IBUF  _2748_ (
    .I(s9_data_i[8]),
    .O(_0236_[8])
  );
IBUF  _2749_ (
    .I(s9_data_i[9]),
    .O(_0236_[9])
  );
OBUF  _2750_ (
    .I(_0237_[0]),
    .O(s9_data_o[0])
  );
OBUF  _2751_ (
    .I(_0237_[1]),
    .O(s9_data_o[1])
  );
OBUF  _2752_ (
    .I(_0237_[10]),
    .O(s9_data_o[10])
  );
OBUF  _2753_ (
    .I(_0237_[11]),
    .O(s9_data_o[11])
  );
OBUF  _2754_ (
    .I(_0237_[12]),
    .O(s9_data_o[12])
  );
OBUF  _2755_ (
    .I(_0237_[13]),
    .O(s9_data_o[13])
  );
OBUF  _2756_ (
    .I(_0237_[14]),
    .O(s9_data_o[14])
  );
OBUF  _2757_ (
    .I(_0237_[15]),
    .O(s9_data_o[15])
  );
OBUF  _2758_ (
    .I(_0237_[16]),
    .O(s9_data_o[16])
  );
OBUF  _2759_ (
    .I(_0237_[17]),
    .O(s9_data_o[17])
  );
OBUF  _2760_ (
    .I(_0237_[18]),
    .O(s9_data_o[18])
  );
OBUF  _2761_ (
    .I(_0237_[19]),
    .O(s9_data_o[19])
  );
OBUF  _2762_ (
    .I(_0237_[2]),
    .O(s9_data_o[2])
  );
OBUF  _2763_ (
    .I(_0237_[20]),
    .O(s9_data_o[20])
  );
OBUF  _2764_ (
    .I(_0237_[21]),
    .O(s9_data_o[21])
  );
OBUF  _2765_ (
    .I(_0237_[22]),
    .O(s9_data_o[22])
  );
OBUF  _2766_ (
    .I(_0237_[23]),
    .O(s9_data_o[23])
  );
OBUF  _2767_ (
    .I(_0237_[24]),
    .O(s9_data_o[24])
  );
OBUF  _2768_ (
    .I(_0237_[25]),
    .O(s9_data_o[25])
  );
OBUF  _2769_ (
    .I(_0237_[26]),
    .O(s9_data_o[26])
  );
OBUF  _2770_ (
    .I(_0237_[27]),
    .O(s9_data_o[27])
  );
OBUF  _2771_ (
    .I(_0237_[28]),
    .O(s9_data_o[28])
  );
OBUF  _2772_ (
    .I(_0237_[29]),
    .O(s9_data_o[29])
  );
OBUF  _2773_ (
    .I(_0237_[3]),
    .O(s9_data_o[3])
  );
OBUF  _2774_ (
    .I(_0237_[30]),
    .O(s9_data_o[30])
  );
OBUF  _2775_ (
    .I(_0237_[31]),
    .O(s9_data_o[31])
  );
OBUF  _2776_ (
    .I(_0237_[4]),
    .O(s9_data_o[4])
  );
OBUF  _2777_ (
    .I(_0237_[5]),
    .O(s9_data_o[5])
  );
OBUF  _2778_ (
    .I(_0237_[6]),
    .O(s9_data_o[6])
  );
OBUF  _2779_ (
    .I(_0237_[7]),
    .O(s9_data_o[7])
  );
OBUF  _2780_ (
    .I(_0237_[8]),
    .O(s9_data_o[8])
  );
OBUF  _2781_ (
    .I(_0237_[9]),
    .O(s9_data_o[9])
  );
IBUF  _2782_ (
    .I(s9_err_i),
    .O(_0238_)
  );
IBUF  _2783_ (
    .I(s9_rty_i),
    .O(_0239_)
  );
OBUF  _2784_ (
    .I(_0240_[0]),
    .O(s9_sel_o[0])
  );
OBUF  _2785_ (
    .I(_0240_[1]),
    .O(s9_sel_o[1])
  );
OBUF  _2786_ (
    .I(_0240_[2]),
    .O(s9_sel_o[2])
  );
OBUF  _2787_ (
    .I(_0240_[3]),
    .O(s9_sel_o[3])
  );
OBUF  _2788_ (
    .I(_0241_),
    .O(s9_stb_o)
  );
OBUF  _2789_ (
    .I(_0242_),
    .O(s9_we_o)
  );
\$paramod$7ef9a024e49224e54bf5d1f376214065d47809cb\wb_conmax_master_if   m0 (
    .clk_i(_0001_),
    .rst_i(_0082_),
    .s0_ack_i(m0s0_ack),
    .s0_addr_o(m0s0_addr),
    .s0_cyc_o(m0s0_cyc),
    .s0_data_i(m0s0_data_i),
    .s0_data_o(m0s0_data_o),
    .s0_err_i(m0s0_err),
    .s0_rty_i(m0s0_rty),
    .s0_sel_o(m0s0_sel),
    .s0_stb_o(m0s0_stb),
    .s0_we_o(m0s0_we),
    .s10_ack_i(m0s10_ack),
    .s10_addr_o(m0s10_addr),
    .s10_cyc_o(m0s10_cyc),
    .s10_data_i(m0s10_data_i),
    .s10_data_o(m0s10_data_o),
    .s10_err_i(m0s10_err),
    .s10_rty_i(m0s10_rty),
    .s10_sel_o(m0s10_sel),
    .s10_stb_o(m0s10_stb),
    .s10_we_o(m0s10_we),
    .s11_ack_i(m0s11_ack),
    .s11_addr_o(m0s11_addr),
    .s11_cyc_o(m0s11_cyc),
    .s11_data_i(m0s11_data_i),
    .s11_data_o(m0s11_data_o),
    .s11_err_i(m0s11_err),
    .s11_rty_i(m0s11_rty),
    .s11_sel_o(m0s11_sel),
    .s11_stb_o(m0s11_stb),
    .s11_we_o(m0s11_we),
    .s12_ack_i(m0s12_ack),
    .s12_addr_o(m0s12_addr),
    .s12_cyc_o(m0s12_cyc),
    .s12_data_i(m0s12_data_i),
    .s12_data_o(m0s12_data_o),
    .s12_err_i(m0s12_err),
    .s12_rty_i(m0s12_rty),
    .s12_sel_o(m0s12_sel),
    .s12_stb_o(m0s12_stb),
    .s12_we_o(m0s12_we),
    .s13_ack_i(m0s13_ack),
    .s13_addr_o(m0s13_addr),
    .s13_cyc_o(m0s13_cyc),
    .s13_data_i(m0s13_data_i),
    .s13_data_o(m0s13_data_o),
    .s13_err_i(m0s13_err),
    .s13_rty_i(m0s13_rty),
    .s13_sel_o(m0s13_sel),
    .s13_stb_o(m0s13_stb),
    .s13_we_o(m0s13_we),
    .s14_ack_i(m0s14_ack),
    .s14_addr_o(m0s14_addr),
    .s14_cyc_o(m0s14_cyc),
    .s14_data_i(m0s14_data_i),
    .s14_data_o(m0s14_data_o),
    .s14_err_i(m0s14_err),
    .s14_rty_i(m0s14_rty),
    .s14_sel_o(m0s14_sel),
    .s14_stb_o(m0s14_stb),
    .s14_we_o(m0s14_we),
    .s15_ack_i(m0s15_ack),
    .s15_addr_o(m0s15_addr),
    .s15_cyc_o(m0s15_cyc),
    .s15_data_i(m0s15_data_i),
    .s15_data_o(m0s15_data_o),
    .s15_err_i(m0s15_err),
    .s15_rty_i(m0s15_rty),
    .s15_sel_o(m0s15_sel),
    .s15_stb_o(m0s15_stb),
    .s15_we_o(m0s15_we),
    .s1_ack_i(m0s1_ack),
    .s1_addr_o(m0s1_addr),
    .s1_cyc_o(m0s1_cyc),
    .s1_data_i(m0s1_data_i),
    .s1_data_o(m0s1_data_o),
    .s1_err_i(m0s1_err),
    .s1_rty_i(m0s1_rty),
    .s1_sel_o(m0s1_sel),
    .s1_stb_o(m0s1_stb),
    .s1_we_o(m0s1_we),
    .s2_ack_i(m0s2_ack),
    .s2_addr_o(m0s2_addr),
    .s2_cyc_o(m0s2_cyc),
    .s2_data_i(m0s2_data_i),
    .s2_data_o(m0s2_data_o),
    .s2_err_i(m0s2_err),
    .s2_rty_i(m0s2_rty),
    .s2_sel_o(m0s2_sel),
    .s2_stb_o(m0s2_stb),
    .s2_we_o(m0s2_we),
    .s3_ack_i(m0s3_ack),
    .s3_addr_o(m0s3_addr),
    .s3_cyc_o(m0s3_cyc),
    .s3_data_i(m0s3_data_i),
    .s3_data_o(m0s3_data_o),
    .s3_err_i(m0s3_err),
    .s3_rty_i(m0s3_rty),
    .s3_sel_o(m0s3_sel),
    .s3_stb_o(m0s3_stb),
    .s3_we_o(m0s3_we),
    .s4_ack_i(m0s4_ack),
    .s4_addr_o(m0s4_addr),
    .s4_cyc_o(m0s4_cyc),
    .s4_data_i(m0s4_data_i),
    .s4_data_o(m0s4_data_o),
    .s4_err_i(m0s4_err),
    .s4_rty_i(m0s4_rty),
    .s4_sel_o(m0s4_sel),
    .s4_stb_o(m0s4_stb),
    .s4_we_o(m0s4_we),
    .s5_ack_i(m0s5_ack),
    .s5_addr_o(m0s5_addr),
    .s5_cyc_o(m0s5_cyc),
    .s5_data_i(m0s5_data_i),
    .s5_data_o(m0s5_data_o),
    .s5_err_i(m0s5_err),
    .s5_rty_i(m0s5_rty),
    .s5_sel_o(m0s5_sel),
    .s5_stb_o(m0s5_stb),
    .s5_we_o(m0s5_we),
    .s6_ack_i(m0s6_ack),
    .s6_addr_o(m0s6_addr),
    .s6_cyc_o(m0s6_cyc),
    .s6_data_i(m0s6_data_i),
    .s6_data_o(m0s6_data_o),
    .s6_err_i(m0s6_err),
    .s6_rty_i(m0s6_rty),
    .s6_sel_o(m0s6_sel),
    .s6_stb_o(m0s6_stb),
    .s6_we_o(m0s6_we),
    .s7_ack_i(m0s7_ack),
    .s7_addr_o(m0s7_addr),
    .s7_cyc_o(m0s7_cyc),
    .s7_data_i(m0s7_data_i),
    .s7_data_o(m0s7_data_o),
    .s7_err_i(m0s7_err),
    .s7_rty_i(m0s7_rty),
    .s7_sel_o(m0s7_sel),
    .s7_stb_o(m0s7_stb),
    .s7_we_o(m0s7_we),
    .s8_ack_i(m0s8_ack),
    .s8_addr_o(m0s8_addr),
    .s8_cyc_o(m0s8_cyc),
    .s8_data_i(m0s8_data_i),
    .s8_data_o(m0s8_data_o),
    .s8_err_i(m0s8_err),
    .s8_rty_i(m0s8_rty),
    .s8_sel_o(m0s8_sel),
    .s8_stb_o(m0s8_stb),
    .s8_we_o(m0s8_we),
    .s9_ack_i(m0s9_ack),
    .s9_addr_o(m0s9_addr),
    .s9_cyc_o(m0s9_cyc),
    .s9_data_i(m0s9_data_i),
    .s9_data_o(m0s9_data_o),
    .s9_err_i(m0s9_err),
    .s9_rty_i(m0s9_rty),
    .s9_sel_o(m0s9_sel),
    .s9_stb_o(m0s9_stb),
    .s9_we_o(m0s9_we),
    .wb_ack_o(_0002_),
    .wb_addr_i(_0003_),
    .wb_cyc_i(_0004_),
    .wb_data_i(_0005_),
    .wb_data_o(_0006_),
    .wb_err_o(_0007_),
    .wb_rty_o(_0008_),
    .wb_sel_i(_0009_),
    .wb_stb_i(_0010_),
    .wb_we_i(_0011_)
  );
\$paramod$7ef9a024e49224e54bf5d1f376214065d47809cb\wb_conmax_master_if   m1 (
    .clk_i(_0001_),
    .rst_i(_0082_),
    .s0_ack_i(m1s0_ack),
    .s0_addr_o(m1s0_addr),
    .s0_cyc_o(m1s0_cyc),
    .s0_data_i(m1s0_data_i),
    .s0_data_o(m1s0_data_o),
    .s0_err_i(m1s0_err),
    .s0_rty_i(m1s0_rty),
    .s0_sel_o(m1s0_sel),
    .s0_stb_o(m1s0_stb),
    .s0_we_o(m1s0_we),
    .s10_ack_i(m1s10_ack),
    .s10_addr_o(m1s10_addr),
    .s10_cyc_o(m1s10_cyc),
    .s10_data_i(m1s10_data_i),
    .s10_data_o(m1s10_data_o),
    .s10_err_i(m1s10_err),
    .s10_rty_i(m1s10_rty),
    .s10_sel_o(m1s10_sel),
    .s10_stb_o(m1s10_stb),
    .s10_we_o(m1s10_we),
    .s11_ack_i(m1s11_ack),
    .s11_addr_o(m1s11_addr),
    .s11_cyc_o(m1s11_cyc),
    .s11_data_i(m1s11_data_i),
    .s11_data_o(m1s11_data_o),
    .s11_err_i(m1s11_err),
    .s11_rty_i(m1s11_rty),
    .s11_sel_o(m1s11_sel),
    .s11_stb_o(m1s11_stb),
    .s11_we_o(m1s11_we),
    .s12_ack_i(m1s12_ack),
    .s12_addr_o(m1s12_addr),
    .s12_cyc_o(m1s12_cyc),
    .s12_data_i(m1s12_data_i),
    .s12_data_o(m1s12_data_o),
    .s12_err_i(m1s12_err),
    .s12_rty_i(m1s12_rty),
    .s12_sel_o(m1s12_sel),
    .s12_stb_o(m1s12_stb),
    .s12_we_o(m1s12_we),
    .s13_ack_i(m1s13_ack),
    .s13_addr_o(m1s13_addr),
    .s13_cyc_o(m1s13_cyc),
    .s13_data_i(m1s13_data_i),
    .s13_data_o(m1s13_data_o),
    .s13_err_i(m1s13_err),
    .s13_rty_i(m1s13_rty),
    .s13_sel_o(m1s13_sel),
    .s13_stb_o(m1s13_stb),
    .s13_we_o(m1s13_we),
    .s14_ack_i(m1s14_ack),
    .s14_addr_o(m1s14_addr),
    .s14_cyc_o(m1s14_cyc),
    .s14_data_i(m1s14_data_i),
    .s14_data_o(m1s14_data_o),
    .s14_err_i(m1s14_err),
    .s14_rty_i(m1s14_rty),
    .s14_sel_o(m1s14_sel),
    .s14_stb_o(m1s14_stb),
    .s14_we_o(m1s14_we),
    .s15_ack_i(m1s15_ack),
    .s15_addr_o(m1s15_addr),
    .s15_cyc_o(m1s15_cyc),
    .s15_data_i(m1s15_data_i),
    .s15_data_o(m1s15_data_o),
    .s15_err_i(m1s15_err),
    .s15_rty_i(m1s15_rty),
    .s15_sel_o(m1s15_sel),
    .s15_stb_o(m1s15_stb),
    .s15_we_o(m1s15_we),
    .s1_ack_i(m1s1_ack),
    .s1_addr_o(m1s1_addr),
    .s1_cyc_o(m1s1_cyc),
    .s1_data_i(m1s1_data_i),
    .s1_data_o(m1s1_data_o),
    .s1_err_i(m1s1_err),
    .s1_rty_i(m1s1_rty),
    .s1_sel_o(m1s1_sel),
    .s1_stb_o(m1s1_stb),
    .s1_we_o(m1s1_we),
    .s2_ack_i(m1s2_ack),
    .s2_addr_o(m1s2_addr),
    .s2_cyc_o(m1s2_cyc),
    .s2_data_i(m1s2_data_i),
    .s2_data_o(m1s2_data_o),
    .s2_err_i(m1s2_err),
    .s2_rty_i(m1s2_rty),
    .s2_sel_o(m1s2_sel),
    .s2_stb_o(m1s2_stb),
    .s2_we_o(m1s2_we),
    .s3_ack_i(m1s3_ack),
    .s3_addr_o(m1s3_addr),
    .s3_cyc_o(m1s3_cyc),
    .s3_data_i(m1s3_data_i),
    .s3_data_o(m1s3_data_o),
    .s3_err_i(m1s3_err),
    .s3_rty_i(m1s3_rty),
    .s3_sel_o(m1s3_sel),
    .s3_stb_o(m1s3_stb),
    .s3_we_o(m1s3_we),
    .s4_ack_i(m1s4_ack),
    .s4_addr_o(m1s4_addr),
    .s4_cyc_o(m1s4_cyc),
    .s4_data_i(m1s4_data_i),
    .s4_data_o(m1s4_data_o),
    .s4_err_i(m1s4_err),
    .s4_rty_i(m1s4_rty),
    .s4_sel_o(m1s4_sel),
    .s4_stb_o(m1s4_stb),
    .s4_we_o(m1s4_we),
    .s5_ack_i(m1s5_ack),
    .s5_addr_o(m1s5_addr),
    .s5_cyc_o(m1s5_cyc),
    .s5_data_i(m1s5_data_i),
    .s5_data_o(m1s5_data_o),
    .s5_err_i(m1s5_err),
    .s5_rty_i(m1s5_rty),
    .s5_sel_o(m1s5_sel),
    .s5_stb_o(m1s5_stb),
    .s5_we_o(m1s5_we),
    .s6_ack_i(m1s6_ack),
    .s6_addr_o(m1s6_addr),
    .s6_cyc_o(m1s6_cyc),
    .s6_data_i(m1s6_data_i),
    .s6_data_o(m1s6_data_o),
    .s6_err_i(m1s6_err),
    .s6_rty_i(m1s6_rty),
    .s6_sel_o(m1s6_sel),
    .s6_stb_o(m1s6_stb),
    .s6_we_o(m1s6_we),
    .s7_ack_i(m1s7_ack),
    .s7_addr_o(m1s7_addr),
    .s7_cyc_o(m1s7_cyc),
    .s7_data_i(m1s7_data_i),
    .s7_data_o(m1s7_data_o),
    .s7_err_i(m1s7_err),
    .s7_rty_i(m1s7_rty),
    .s7_sel_o(m1s7_sel),
    .s7_stb_o(m1s7_stb),
    .s7_we_o(m1s7_we),
    .s8_ack_i(m1s8_ack),
    .s8_addr_o(m1s8_addr),
    .s8_cyc_o(m1s8_cyc),
    .s8_data_i(m1s8_data_i),
    .s8_data_o(m1s8_data_o),
    .s8_err_i(m1s8_err),
    .s8_rty_i(m1s8_rty),
    .s8_sel_o(m1s8_sel),
    .s8_stb_o(m1s8_stb),
    .s8_we_o(m1s8_we),
    .s9_ack_i(m1s9_ack),
    .s9_addr_o(m1s9_addr),
    .s9_cyc_o(m1s9_cyc),
    .s9_data_i(m1s9_data_i),
    .s9_data_o(m1s9_data_o),
    .s9_err_i(m1s9_err),
    .s9_rty_i(m1s9_rty),
    .s9_sel_o(m1s9_sel),
    .s9_stb_o(m1s9_stb),
    .s9_we_o(m1s9_we),
    .wb_ack_o(_0012_),
    .wb_addr_i(_0013_),
    .wb_cyc_i(_0014_),
    .wb_data_i(_0015_),
    .wb_data_o(_0016_),
    .wb_err_o(_0017_),
    .wb_rty_o(_0018_),
    .wb_sel_i(_0019_),
    .wb_stb_i(_0020_),
    .wb_we_i(_0021_)
  );
\$paramod$7ef9a024e49224e54bf5d1f376214065d47809cb\wb_conmax_master_if   m2 (
    .clk_i(_0001_),
    .rst_i(_0082_),
    .s0_ack_i(m2s0_ack),
    .s0_addr_o(m2s0_addr),
    .s0_cyc_o(m2s0_cyc),
    .s0_data_i(m2s0_data_i),
    .s0_data_o(m2s0_data_o),
    .s0_err_i(m2s0_err),
    .s0_rty_i(m2s0_rty),
    .s0_sel_o(m2s0_sel),
    .s0_stb_o(m2s0_stb),
    .s0_we_o(m2s0_we),
    .s10_ack_i(m2s10_ack),
    .s10_addr_o(m2s10_addr),
    .s10_cyc_o(m2s10_cyc),
    .s10_data_i(m2s10_data_i),
    .s10_data_o(m2s10_data_o),
    .s10_err_i(m2s10_err),
    .s10_rty_i(m2s10_rty),
    .s10_sel_o(m2s10_sel),
    .s10_stb_o(m2s10_stb),
    .s10_we_o(m2s10_we),
    .s11_ack_i(m2s11_ack),
    .s11_addr_o(m2s11_addr),
    .s11_cyc_o(m2s11_cyc),
    .s11_data_i(m2s11_data_i),
    .s11_data_o(m2s11_data_o),
    .s11_err_i(m2s11_err),
    .s11_rty_i(m2s11_rty),
    .s11_sel_o(m2s11_sel),
    .s11_stb_o(m2s11_stb),
    .s11_we_o(m2s11_we),
    .s12_ack_i(m2s12_ack),
    .s12_addr_o(m2s12_addr),
    .s12_cyc_o(m2s12_cyc),
    .s12_data_i(m2s12_data_i),
    .s12_data_o(m2s12_data_o),
    .s12_err_i(m2s12_err),
    .s12_rty_i(m2s12_rty),
    .s12_sel_o(m2s12_sel),
    .s12_stb_o(m2s12_stb),
    .s12_we_o(m2s12_we),
    .s13_ack_i(m2s13_ack),
    .s13_addr_o(m2s13_addr),
    .s13_cyc_o(m2s13_cyc),
    .s13_data_i(m2s13_data_i),
    .s13_data_o(m2s13_data_o),
    .s13_err_i(m2s13_err),
    .s13_rty_i(m2s13_rty),
    .s13_sel_o(m2s13_sel),
    .s13_stb_o(m2s13_stb),
    .s13_we_o(m2s13_we),
    .s14_ack_i(m2s14_ack),
    .s14_addr_o(m2s14_addr),
    .s14_cyc_o(m2s14_cyc),
    .s14_data_i(m2s14_data_i),
    .s14_data_o(m2s14_data_o),
    .s14_err_i(m2s14_err),
    .s14_rty_i(m2s14_rty),
    .s14_sel_o(m2s14_sel),
    .s14_stb_o(m2s14_stb),
    .s14_we_o(m2s14_we),
    .s15_ack_i(m2s15_ack),
    .s15_addr_o(m2s15_addr),
    .s15_cyc_o(m2s15_cyc),
    .s15_data_i(m2s15_data_i),
    .s15_data_o(m2s15_data_o),
    .s15_err_i(m2s15_err),
    .s15_rty_i(m2s15_rty),
    .s15_sel_o(m2s15_sel),
    .s15_stb_o(m2s15_stb),
    .s15_we_o(m2s15_we),
    .s1_ack_i(m2s1_ack),
    .s1_addr_o(m2s1_addr),
    .s1_cyc_o(m2s1_cyc),
    .s1_data_i(m2s1_data_i),
    .s1_data_o(m2s1_data_o),
    .s1_err_i(m2s1_err),
    .s1_rty_i(m2s1_rty),
    .s1_sel_o(m2s1_sel),
    .s1_stb_o(m2s1_stb),
    .s1_we_o(m2s1_we),
    .s2_ack_i(m2s2_ack),
    .s2_addr_o(m2s2_addr),
    .s2_cyc_o(m2s2_cyc),
    .s2_data_i(m2s2_data_i),
    .s2_data_o(m2s2_data_o),
    .s2_err_i(m2s2_err),
    .s2_rty_i(m2s2_rty),
    .s2_sel_o(m2s2_sel),
    .s2_stb_o(m2s2_stb),
    .s2_we_o(m2s2_we),
    .s3_ack_i(m2s3_ack),
    .s3_addr_o(m2s3_addr),
    .s3_cyc_o(m2s3_cyc),
    .s3_data_i(m2s3_data_i),
    .s3_data_o(m2s3_data_o),
    .s3_err_i(m2s3_err),
    .s3_rty_i(m2s3_rty),
    .s3_sel_o(m2s3_sel),
    .s3_stb_o(m2s3_stb),
    .s3_we_o(m2s3_we),
    .s4_ack_i(m2s4_ack),
    .s4_addr_o(m2s4_addr),
    .s4_cyc_o(m2s4_cyc),
    .s4_data_i(m2s4_data_i),
    .s4_data_o(m2s4_data_o),
    .s4_err_i(m2s4_err),
    .s4_rty_i(m2s4_rty),
    .s4_sel_o(m2s4_sel),
    .s4_stb_o(m2s4_stb),
    .s4_we_o(m2s4_we),
    .s5_ack_i(m2s5_ack),
    .s5_addr_o(m2s5_addr),
    .s5_cyc_o(m2s5_cyc),
    .s5_data_i(m2s5_data_i),
    .s5_data_o(m2s5_data_o),
    .s5_err_i(m2s5_err),
    .s5_rty_i(m2s5_rty),
    .s5_sel_o(m2s5_sel),
    .s5_stb_o(m2s5_stb),
    .s5_we_o(m2s5_we),
    .s6_ack_i(m2s6_ack),
    .s6_addr_o(m2s6_addr),
    .s6_cyc_o(m2s6_cyc),
    .s6_data_i(m2s6_data_i),
    .s6_data_o(m2s6_data_o),
    .s6_err_i(m2s6_err),
    .s6_rty_i(m2s6_rty),
    .s6_sel_o(m2s6_sel),
    .s6_stb_o(m2s6_stb),
    .s6_we_o(m2s6_we),
    .s7_ack_i(m2s7_ack),
    .s7_addr_o(m2s7_addr),
    .s7_cyc_o(m2s7_cyc),
    .s7_data_i(m2s7_data_i),
    .s7_data_o(m2s7_data_o),
    .s7_err_i(m2s7_err),
    .s7_rty_i(m2s7_rty),
    .s7_sel_o(m2s7_sel),
    .s7_stb_o(m2s7_stb),
    .s7_we_o(m2s7_we),
    .s8_ack_i(m2s8_ack),
    .s8_addr_o(m2s8_addr),
    .s8_cyc_o(m2s8_cyc),
    .s8_data_i(m2s8_data_i),
    .s8_data_o(m2s8_data_o),
    .s8_err_i(m2s8_err),
    .s8_rty_i(m2s8_rty),
    .s8_sel_o(m2s8_sel),
    .s8_stb_o(m2s8_stb),
    .s8_we_o(m2s8_we),
    .s9_ack_i(m2s9_ack),
    .s9_addr_o(m2s9_addr),
    .s9_cyc_o(m2s9_cyc),
    .s9_data_i(m2s9_data_i),
    .s9_data_o(m2s9_data_o),
    .s9_err_i(m2s9_err),
    .s9_rty_i(m2s9_rty),
    .s9_sel_o(m2s9_sel),
    .s9_stb_o(m2s9_stb),
    .s9_we_o(m2s9_we),
    .wb_ack_o(_0022_),
    .wb_addr_i(_0023_),
    .wb_cyc_i(_0024_),
    .wb_data_i(_0025_),
    .wb_data_o(_0026_),
    .wb_err_o(_0027_),
    .wb_rty_o(_0028_),
    .wb_sel_i(_0029_),
    .wb_stb_i(_0030_),
    .wb_we_i(_0031_)
  );
\$paramod$7ef9a024e49224e54bf5d1f376214065d47809cb\wb_conmax_master_if   m3 (
    .clk_i(_0001_),
    .rst_i(_0082_),
    .s0_ack_i(m3s0_ack),
    .s0_addr_o(m3s0_addr),
    .s0_cyc_o(m3s0_cyc),
    .s0_data_i(m3s0_data_i),
    .s0_data_o(m3s0_data_o),
    .s0_err_i(m3s0_err),
    .s0_rty_i(m3s0_rty),
    .s0_sel_o(m3s0_sel),
    .s0_stb_o(m3s0_stb),
    .s0_we_o(m3s0_we),
    .s10_ack_i(m3s10_ack),
    .s10_addr_o(m3s10_addr),
    .s10_cyc_o(m3s10_cyc),
    .s10_data_i(m3s10_data_i),
    .s10_data_o(m3s10_data_o),
    .s10_err_i(m3s10_err),
    .s10_rty_i(m3s10_rty),
    .s10_sel_o(m3s10_sel),
    .s10_stb_o(m3s10_stb),
    .s10_we_o(m3s10_we),
    .s11_ack_i(m3s11_ack),
    .s11_addr_o(m3s11_addr),
    .s11_cyc_o(m3s11_cyc),
    .s11_data_i(m3s11_data_i),
    .s11_data_o(m3s11_data_o),
    .s11_err_i(m3s11_err),
    .s11_rty_i(m3s11_rty),
    .s11_sel_o(m3s11_sel),
    .s11_stb_o(m3s11_stb),
    .s11_we_o(m3s11_we),
    .s12_ack_i(m3s12_ack),
    .s12_addr_o(m3s12_addr),
    .s12_cyc_o(m3s12_cyc),
    .s12_data_i(m3s12_data_i),
    .s12_data_o(m3s12_data_o),
    .s12_err_i(m3s12_err),
    .s12_rty_i(m3s12_rty),
    .s12_sel_o(m3s12_sel),
    .s12_stb_o(m3s12_stb),
    .s12_we_o(m3s12_we),
    .s13_ack_i(m3s13_ack),
    .s13_addr_o(m3s13_addr),
    .s13_cyc_o(m3s13_cyc),
    .s13_data_i(m3s13_data_i),
    .s13_data_o(m3s13_data_o),
    .s13_err_i(m3s13_err),
    .s13_rty_i(m3s13_rty),
    .s13_sel_o(m3s13_sel),
    .s13_stb_o(m3s13_stb),
    .s13_we_o(m3s13_we),
    .s14_ack_i(m3s14_ack),
    .s14_addr_o(m3s14_addr),
    .s14_cyc_o(m3s14_cyc),
    .s14_data_i(m3s14_data_i),
    .s14_data_o(m3s14_data_o),
    .s14_err_i(m3s14_err),
    .s14_rty_i(m3s14_rty),
    .s14_sel_o(m3s14_sel),
    .s14_stb_o(m3s14_stb),
    .s14_we_o(m3s14_we),
    .s15_ack_i(m3s15_ack),
    .s15_addr_o(m3s15_addr),
    .s15_cyc_o(m3s15_cyc),
    .s15_data_i(m3s15_data_i),
    .s15_data_o(m3s15_data_o),
    .s15_err_i(m3s15_err),
    .s15_rty_i(m3s15_rty),
    .s15_sel_o(m3s15_sel),
    .s15_stb_o(m3s15_stb),
    .s15_we_o(m3s15_we),
    .s1_ack_i(m3s1_ack),
    .s1_addr_o(m3s1_addr),
    .s1_cyc_o(m3s1_cyc),
    .s1_data_i(m3s1_data_i),
    .s1_data_o(m3s1_data_o),
    .s1_err_i(m3s1_err),
    .s1_rty_i(m3s1_rty),
    .s1_sel_o(m3s1_sel),
    .s1_stb_o(m3s1_stb),
    .s1_we_o(m3s1_we),
    .s2_ack_i(m3s2_ack),
    .s2_addr_o(m3s2_addr),
    .s2_cyc_o(m3s2_cyc),
    .s2_data_i(m3s2_data_i),
    .s2_data_o(m3s2_data_o),
    .s2_err_i(m3s2_err),
    .s2_rty_i(m3s2_rty),
    .s2_sel_o(m3s2_sel),
    .s2_stb_o(m3s2_stb),
    .s2_we_o(m3s2_we),
    .s3_ack_i(m3s3_ack),
    .s3_addr_o(m3s3_addr),
    .s3_cyc_o(m3s3_cyc),
    .s3_data_i(m3s3_data_i),
    .s3_data_o(m3s3_data_o),
    .s3_err_i(m3s3_err),
    .s3_rty_i(m3s3_rty),
    .s3_sel_o(m3s3_sel),
    .s3_stb_o(m3s3_stb),
    .s3_we_o(m3s3_we),
    .s4_ack_i(m3s4_ack),
    .s4_addr_o(m3s4_addr),
    .s4_cyc_o(m3s4_cyc),
    .s4_data_i(m3s4_data_i),
    .s4_data_o(m3s4_data_o),
    .s4_err_i(m3s4_err),
    .s4_rty_i(m3s4_rty),
    .s4_sel_o(m3s4_sel),
    .s4_stb_o(m3s4_stb),
    .s4_we_o(m3s4_we),
    .s5_ack_i(m3s5_ack),
    .s5_addr_o(m3s5_addr),
    .s5_cyc_o(m3s5_cyc),
    .s5_data_i(m3s5_data_i),
    .s5_data_o(m3s5_data_o),
    .s5_err_i(m3s5_err),
    .s5_rty_i(m3s5_rty),
    .s5_sel_o(m3s5_sel),
    .s5_stb_o(m3s5_stb),
    .s5_we_o(m3s5_we),
    .s6_ack_i(m3s6_ack),
    .s6_addr_o(m3s6_addr),
    .s6_cyc_o(m3s6_cyc),
    .s6_data_i(m3s6_data_i),
    .s6_data_o(m3s6_data_o),
    .s6_err_i(m3s6_err),
    .s6_rty_i(m3s6_rty),
    .s6_sel_o(m3s6_sel),
    .s6_stb_o(m3s6_stb),
    .s6_we_o(m3s6_we),
    .s7_ack_i(m3s7_ack),
    .s7_addr_o(m3s7_addr),
    .s7_cyc_o(m3s7_cyc),
    .s7_data_i(m3s7_data_i),
    .s7_data_o(m3s7_data_o),
    .s7_err_i(m3s7_err),
    .s7_rty_i(m3s7_rty),
    .s7_sel_o(m3s7_sel),
    .s7_stb_o(m3s7_stb),
    .s7_we_o(m3s7_we),
    .s8_ack_i(m3s8_ack),
    .s8_addr_o(m3s8_addr),
    .s8_cyc_o(m3s8_cyc),
    .s8_data_i(m3s8_data_i),
    .s8_data_o(m3s8_data_o),
    .s8_err_i(m3s8_err),
    .s8_rty_i(m3s8_rty),
    .s8_sel_o(m3s8_sel),
    .s8_stb_o(m3s8_stb),
    .s8_we_o(m3s8_we),
    .s9_ack_i(m3s9_ack),
    .s9_addr_o(m3s9_addr),
    .s9_cyc_o(m3s9_cyc),
    .s9_data_i(m3s9_data_i),
    .s9_data_o(m3s9_data_o),
    .s9_err_i(m3s9_err),
    .s9_rty_i(m3s9_rty),
    .s9_sel_o(m3s9_sel),
    .s9_stb_o(m3s9_stb),
    .s9_we_o(m3s9_we),
    .wb_ack_o(_0032_),
    .wb_addr_i(_0033_),
    .wb_cyc_i(_0034_),
    .wb_data_i(_0035_),
    .wb_data_o(_0036_),
    .wb_err_o(_0037_),
    .wb_rty_o(_0038_),
    .wb_sel_i(_0039_),
    .wb_stb_i(_0040_),
    .wb_we_i(_0041_)
  );
\$paramod$7ef9a024e49224e54bf5d1f376214065d47809cb\wb_conmax_master_if   m4 (
    .clk_i(_0001_),
    .rst_i(_0082_),
    .s0_ack_i(m4s0_ack),
    .s0_addr_o(m4s0_addr),
    .s0_cyc_o(m4s0_cyc),
    .s0_data_i(m4s0_data_i),
    .s0_data_o(m4s0_data_o),
    .s0_err_i(m4s0_err),
    .s0_rty_i(m4s0_rty),
    .s0_sel_o(m4s0_sel),
    .s0_stb_o(m4s0_stb),
    .s0_we_o(m4s0_we),
    .s10_ack_i(m4s10_ack),
    .s10_addr_o(m4s10_addr),
    .s10_cyc_o(m4s10_cyc),
    .s10_data_i(m4s10_data_i),
    .s10_data_o(m4s10_data_o),
    .s10_err_i(m4s10_err),
    .s10_rty_i(m4s10_rty),
    .s10_sel_o(m4s10_sel),
    .s10_stb_o(m4s10_stb),
    .s10_we_o(m4s10_we),
    .s11_ack_i(m4s11_ack),
    .s11_addr_o(m4s11_addr),
    .s11_cyc_o(m4s11_cyc),
    .s11_data_i(m4s11_data_i),
    .s11_data_o(m4s11_data_o),
    .s11_err_i(m4s11_err),
    .s11_rty_i(m4s11_rty),
    .s11_sel_o(m4s11_sel),
    .s11_stb_o(m4s11_stb),
    .s11_we_o(m4s11_we),
    .s12_ack_i(m4s12_ack),
    .s12_addr_o(m4s12_addr),
    .s12_cyc_o(m4s12_cyc),
    .s12_data_i(m4s12_data_i),
    .s12_data_o(m4s12_data_o),
    .s12_err_i(m4s12_err),
    .s12_rty_i(m4s12_rty),
    .s12_sel_o(m4s12_sel),
    .s12_stb_o(m4s12_stb),
    .s12_we_o(m4s12_we),
    .s13_ack_i(m4s13_ack),
    .s13_addr_o(m4s13_addr),
    .s13_cyc_o(m4s13_cyc),
    .s13_data_i(m4s13_data_i),
    .s13_data_o(m4s13_data_o),
    .s13_err_i(m4s13_err),
    .s13_rty_i(m4s13_rty),
    .s13_sel_o(m4s13_sel),
    .s13_stb_o(m4s13_stb),
    .s13_we_o(m4s13_we),
    .s14_ack_i(m4s14_ack),
    .s14_addr_o(m4s14_addr),
    .s14_cyc_o(m4s14_cyc),
    .s14_data_i(m4s14_data_i),
    .s14_data_o(m4s14_data_o),
    .s14_err_i(m4s14_err),
    .s14_rty_i(m4s14_rty),
    .s14_sel_o(m4s14_sel),
    .s14_stb_o(m4s14_stb),
    .s14_we_o(m4s14_we),
    .s15_ack_i(m4s15_ack),
    .s15_addr_o(m4s15_addr),
    .s15_cyc_o(m4s15_cyc),
    .s15_data_i(m4s15_data_i),
    .s15_data_o(m4s15_data_o),
    .s15_err_i(m4s15_err),
    .s15_rty_i(m4s15_rty),
    .s15_sel_o(m4s15_sel),
    .s15_stb_o(m4s15_stb),
    .s15_we_o(m4s15_we),
    .s1_ack_i(m4s1_ack),
    .s1_addr_o(m4s1_addr),
    .s1_cyc_o(m4s1_cyc),
    .s1_data_i(m4s1_data_i),
    .s1_data_o(m4s1_data_o),
    .s1_err_i(m4s1_err),
    .s1_rty_i(m4s1_rty),
    .s1_sel_o(m4s1_sel),
    .s1_stb_o(m4s1_stb),
    .s1_we_o(m4s1_we),
    .s2_ack_i(m4s2_ack),
    .s2_addr_o(m4s2_addr),
    .s2_cyc_o(m4s2_cyc),
    .s2_data_i(m4s2_data_i),
    .s2_data_o(m4s2_data_o),
    .s2_err_i(m4s2_err),
    .s2_rty_i(m4s2_rty),
    .s2_sel_o(m4s2_sel),
    .s2_stb_o(m4s2_stb),
    .s2_we_o(m4s2_we),
    .s3_ack_i(m4s3_ack),
    .s3_addr_o(m4s3_addr),
    .s3_cyc_o(m4s3_cyc),
    .s3_data_i(m4s3_data_i),
    .s3_data_o(m4s3_data_o),
    .s3_err_i(m4s3_err),
    .s3_rty_i(m4s3_rty),
    .s3_sel_o(m4s3_sel),
    .s3_stb_o(m4s3_stb),
    .s3_we_o(m4s3_we),
    .s4_ack_i(m4s4_ack),
    .s4_addr_o(m4s4_addr),
    .s4_cyc_o(m4s4_cyc),
    .s4_data_i(m4s4_data_i),
    .s4_data_o(m4s4_data_o),
    .s4_err_i(m4s4_err),
    .s4_rty_i(m4s4_rty),
    .s4_sel_o(m4s4_sel),
    .s4_stb_o(m4s4_stb),
    .s4_we_o(m4s4_we),
    .s5_ack_i(m4s5_ack),
    .s5_addr_o(m4s5_addr),
    .s5_cyc_o(m4s5_cyc),
    .s5_data_i(m4s5_data_i),
    .s5_data_o(m4s5_data_o),
    .s5_err_i(m4s5_err),
    .s5_rty_i(m4s5_rty),
    .s5_sel_o(m4s5_sel),
    .s5_stb_o(m4s5_stb),
    .s5_we_o(m4s5_we),
    .s6_ack_i(m4s6_ack),
    .s6_addr_o(m4s6_addr),
    .s6_cyc_o(m4s6_cyc),
    .s6_data_i(m4s6_data_i),
    .s6_data_o(m4s6_data_o),
    .s6_err_i(m4s6_err),
    .s6_rty_i(m4s6_rty),
    .s6_sel_o(m4s6_sel),
    .s6_stb_o(m4s6_stb),
    .s6_we_o(m4s6_we),
    .s7_ack_i(m4s7_ack),
    .s7_addr_o(m4s7_addr),
    .s7_cyc_o(m4s7_cyc),
    .s7_data_i(m4s7_data_i),
    .s7_data_o(m4s7_data_o),
    .s7_err_i(m4s7_err),
    .s7_rty_i(m4s7_rty),
    .s7_sel_o(m4s7_sel),
    .s7_stb_o(m4s7_stb),
    .s7_we_o(m4s7_we),
    .s8_ack_i(m4s8_ack),
    .s8_addr_o(m4s8_addr),
    .s8_cyc_o(m4s8_cyc),
    .s8_data_i(m4s8_data_i),
    .s8_data_o(m4s8_data_o),
    .s8_err_i(m4s8_err),
    .s8_rty_i(m4s8_rty),
    .s8_sel_o(m4s8_sel),
    .s8_stb_o(m4s8_stb),
    .s8_we_o(m4s8_we),
    .s9_ack_i(m4s9_ack),
    .s9_addr_o(m4s9_addr),
    .s9_cyc_o(m4s9_cyc),
    .s9_data_i(m4s9_data_i),
    .s9_data_o(m4s9_data_o),
    .s9_err_i(m4s9_err),
    .s9_rty_i(m4s9_rty),
    .s9_sel_o(m4s9_sel),
    .s9_stb_o(m4s9_stb),
    .s9_we_o(m4s9_we),
    .wb_ack_o(_0042_),
    .wb_addr_i(_0043_),
    .wb_cyc_i(_0044_),
    .wb_data_i(_0045_),
    .wb_data_o(_0046_),
    .wb_err_o(_0047_),
    .wb_rty_o(_0048_),
    .wb_sel_i(_0049_),
    .wb_stb_i(_0050_),
    .wb_we_i(_0051_)
  );
\$paramod$7ef9a024e49224e54bf5d1f376214065d47809cb\wb_conmax_master_if   m5 (
    .clk_i(_0001_),
    .rst_i(_0082_),
    .s0_ack_i(m5s0_ack),
    .s0_addr_o(m5s0_addr),
    .s0_cyc_o(m5s0_cyc),
    .s0_data_i(m5s0_data_i),
    .s0_data_o(m5s0_data_o),
    .s0_err_i(m5s0_err),
    .s0_rty_i(m5s0_rty),
    .s0_sel_o(m5s0_sel),
    .s0_stb_o(m5s0_stb),
    .s0_we_o(m5s0_we),
    .s10_ack_i(m5s10_ack),
    .s10_addr_o(m5s10_addr),
    .s10_cyc_o(m5s10_cyc),
    .s10_data_i(m5s10_data_i),
    .s10_data_o(m5s10_data_o),
    .s10_err_i(m5s10_err),
    .s10_rty_i(m5s10_rty),
    .s10_sel_o(m5s10_sel),
    .s10_stb_o(m5s10_stb),
    .s10_we_o(m5s10_we),
    .s11_ack_i(m5s11_ack),
    .s11_addr_o(m5s11_addr),
    .s11_cyc_o(m5s11_cyc),
    .s11_data_i(m5s11_data_i),
    .s11_data_o(m5s11_data_o),
    .s11_err_i(m5s11_err),
    .s11_rty_i(m5s11_rty),
    .s11_sel_o(m5s11_sel),
    .s11_stb_o(m5s11_stb),
    .s11_we_o(m5s11_we),
    .s12_ack_i(m5s12_ack),
    .s12_addr_o(m5s12_addr),
    .s12_cyc_o(m5s12_cyc),
    .s12_data_i(m5s12_data_i),
    .s12_data_o(m5s12_data_o),
    .s12_err_i(m5s12_err),
    .s12_rty_i(m5s12_rty),
    .s12_sel_o(m5s12_sel),
    .s12_stb_o(m5s12_stb),
    .s12_we_o(m5s12_we),
    .s13_ack_i(m5s13_ack),
    .s13_addr_o(m5s13_addr),
    .s13_cyc_o(m5s13_cyc),
    .s13_data_i(m5s13_data_i),
    .s13_data_o(m5s13_data_o),
    .s13_err_i(m5s13_err),
    .s13_rty_i(m5s13_rty),
    .s13_sel_o(m5s13_sel),
    .s13_stb_o(m5s13_stb),
    .s13_we_o(m5s13_we),
    .s14_ack_i(m5s14_ack),
    .s14_addr_o(m5s14_addr),
    .s14_cyc_o(m5s14_cyc),
    .s14_data_i(m5s14_data_i),
    .s14_data_o(m5s14_data_o),
    .s14_err_i(m5s14_err),
    .s14_rty_i(m5s14_rty),
    .s14_sel_o(m5s14_sel),
    .s14_stb_o(m5s14_stb),
    .s14_we_o(m5s14_we),
    .s15_ack_i(m5s15_ack),
    .s15_addr_o(m5s15_addr),
    .s15_cyc_o(m5s15_cyc),
    .s15_data_i(m5s15_data_i),
    .s15_data_o(m5s15_data_o),
    .s15_err_i(m5s15_err),
    .s15_rty_i(m5s15_rty),
    .s15_sel_o(m5s15_sel),
    .s15_stb_o(m5s15_stb),
    .s15_we_o(m5s15_we),
    .s1_ack_i(m5s1_ack),
    .s1_addr_o(m5s1_addr),
    .s1_cyc_o(m5s1_cyc),
    .s1_data_i(m5s1_data_i),
    .s1_data_o(m5s1_data_o),
    .s1_err_i(m5s1_err),
    .s1_rty_i(m5s1_rty),
    .s1_sel_o(m5s1_sel),
    .s1_stb_o(m5s1_stb),
    .s1_we_o(m5s1_we),
    .s2_ack_i(m5s2_ack),
    .s2_addr_o(m5s2_addr),
    .s2_cyc_o(m5s2_cyc),
    .s2_data_i(m5s2_data_i),
    .s2_data_o(m5s2_data_o),
    .s2_err_i(m5s2_err),
    .s2_rty_i(m5s2_rty),
    .s2_sel_o(m5s2_sel),
    .s2_stb_o(m5s2_stb),
    .s2_we_o(m5s2_we),
    .s3_ack_i(m5s3_ack),
    .s3_addr_o(m5s3_addr),
    .s3_cyc_o(m5s3_cyc),
    .s3_data_i(m5s3_data_i),
    .s3_data_o(m5s3_data_o),
    .s3_err_i(m5s3_err),
    .s3_rty_i(m5s3_rty),
    .s3_sel_o(m5s3_sel),
    .s3_stb_o(m5s3_stb),
    .s3_we_o(m5s3_we),
    .s4_ack_i(m5s4_ack),
    .s4_addr_o(m5s4_addr),
    .s4_cyc_o(m5s4_cyc),
    .s4_data_i(m5s4_data_i),
    .s4_data_o(m5s4_data_o),
    .s4_err_i(m5s4_err),
    .s4_rty_i(m5s4_rty),
    .s4_sel_o(m5s4_sel),
    .s4_stb_o(m5s4_stb),
    .s4_we_o(m5s4_we),
    .s5_ack_i(m5s5_ack),
    .s5_addr_o(m5s5_addr),
    .s5_cyc_o(m5s5_cyc),
    .s5_data_i(m5s5_data_i),
    .s5_data_o(m5s5_data_o),
    .s5_err_i(m5s5_err),
    .s5_rty_i(m5s5_rty),
    .s5_sel_o(m5s5_sel),
    .s5_stb_o(m5s5_stb),
    .s5_we_o(m5s5_we),
    .s6_ack_i(m5s6_ack),
    .s6_addr_o(m5s6_addr),
    .s6_cyc_o(m5s6_cyc),
    .s6_data_i(m5s6_data_i),
    .s6_data_o(m5s6_data_o),
    .s6_err_i(m5s6_err),
    .s6_rty_i(m5s6_rty),
    .s6_sel_o(m5s6_sel),
    .s6_stb_o(m5s6_stb),
    .s6_we_o(m5s6_we),
    .s7_ack_i(m5s7_ack),
    .s7_addr_o(m5s7_addr),
    .s7_cyc_o(m5s7_cyc),
    .s7_data_i(m5s7_data_i),
    .s7_data_o(m5s7_data_o),
    .s7_err_i(m5s7_err),
    .s7_rty_i(m5s7_rty),
    .s7_sel_o(m5s7_sel),
    .s7_stb_o(m5s7_stb),
    .s7_we_o(m5s7_we),
    .s8_ack_i(m5s8_ack),
    .s8_addr_o(m5s8_addr),
    .s8_cyc_o(m5s8_cyc),
    .s8_data_i(m5s8_data_i),
    .s8_data_o(m5s8_data_o),
    .s8_err_i(m5s8_err),
    .s8_rty_i(m5s8_rty),
    .s8_sel_o(m5s8_sel),
    .s8_stb_o(m5s8_stb),
    .s8_we_o(m5s8_we),
    .s9_ack_i(m5s9_ack),
    .s9_addr_o(m5s9_addr),
    .s9_cyc_o(m5s9_cyc),
    .s9_data_i(m5s9_data_i),
    .s9_data_o(m5s9_data_o),
    .s9_err_i(m5s9_err),
    .s9_rty_i(m5s9_rty),
    .s9_sel_o(m5s9_sel),
    .s9_stb_o(m5s9_stb),
    .s9_we_o(m5s9_we),
    .wb_ack_o(_0052_),
    .wb_addr_i(_0053_),
    .wb_cyc_i(_0054_),
    .wb_data_i(_0055_),
    .wb_data_o(_0056_),
    .wb_err_o(_0057_),
    .wb_rty_o(_0058_),
    .wb_sel_i(_0059_),
    .wb_stb_i(_0060_),
    .wb_we_i(_0061_)
  );
\$paramod$7ef9a024e49224e54bf5d1f376214065d47809cb\wb_conmax_master_if   m6 (
    .clk_i(_0001_),
    .rst_i(_0082_),
    .s0_ack_i(m6s0_ack),
    .s0_addr_o(m6s0_addr),
    .s0_cyc_o(m6s0_cyc),
    .s0_data_i(m6s0_data_i),
    .s0_data_o(m6s0_data_o),
    .s0_err_i(m6s0_err),
    .s0_rty_i(m6s0_rty),
    .s0_sel_o(m6s0_sel),
    .s0_stb_o(m6s0_stb),
    .s0_we_o(m6s0_we),
    .s10_ack_i(m6s10_ack),
    .s10_addr_o(m6s10_addr),
    .s10_cyc_o(m6s10_cyc),
    .s10_data_i(m6s10_data_i),
    .s10_data_o(m6s10_data_o),
    .s10_err_i(m6s10_err),
    .s10_rty_i(m6s10_rty),
    .s10_sel_o(m6s10_sel),
    .s10_stb_o(m6s10_stb),
    .s10_we_o(m6s10_we),
    .s11_ack_i(m6s11_ack),
    .s11_addr_o(m6s11_addr),
    .s11_cyc_o(m6s11_cyc),
    .s11_data_i(m6s11_data_i),
    .s11_data_o(m6s11_data_o),
    .s11_err_i(m6s11_err),
    .s11_rty_i(m6s11_rty),
    .s11_sel_o(m6s11_sel),
    .s11_stb_o(m6s11_stb),
    .s11_we_o(m6s11_we),
    .s12_ack_i(m6s12_ack),
    .s12_addr_o(m6s12_addr),
    .s12_cyc_o(m6s12_cyc),
    .s12_data_i(m6s12_data_i),
    .s12_data_o(m6s12_data_o),
    .s12_err_i(m6s12_err),
    .s12_rty_i(m6s12_rty),
    .s12_sel_o(m6s12_sel),
    .s12_stb_o(m6s12_stb),
    .s12_we_o(m6s12_we),
    .s13_ack_i(m6s13_ack),
    .s13_addr_o(m6s13_addr),
    .s13_cyc_o(m6s13_cyc),
    .s13_data_i(m6s13_data_i),
    .s13_data_o(m6s13_data_o),
    .s13_err_i(m6s13_err),
    .s13_rty_i(m6s13_rty),
    .s13_sel_o(m6s13_sel),
    .s13_stb_o(m6s13_stb),
    .s13_we_o(m6s13_we),
    .s14_ack_i(m6s14_ack),
    .s14_addr_o(m6s14_addr),
    .s14_cyc_o(m6s14_cyc),
    .s14_data_i(m6s14_data_i),
    .s14_data_o(m6s14_data_o),
    .s14_err_i(m6s14_err),
    .s14_rty_i(m6s14_rty),
    .s14_sel_o(m6s14_sel),
    .s14_stb_o(m6s14_stb),
    .s14_we_o(m6s14_we),
    .s15_ack_i(m6s15_ack),
    .s15_addr_o(m6s15_addr),
    .s15_cyc_o(m6s15_cyc),
    .s15_data_i(m6s15_data_i),
    .s15_data_o(m6s15_data_o),
    .s15_err_i(m6s15_err),
    .s15_rty_i(m6s15_rty),
    .s15_sel_o(m6s15_sel),
    .s15_stb_o(m6s15_stb),
    .s15_we_o(m6s15_we),
    .s1_ack_i(m6s1_ack),
    .s1_addr_o(m6s1_addr),
    .s1_cyc_o(m6s1_cyc),
    .s1_data_i(m6s1_data_i),
    .s1_data_o(m6s1_data_o),
    .s1_err_i(m6s1_err),
    .s1_rty_i(m6s1_rty),
    .s1_sel_o(m6s1_sel),
    .s1_stb_o(m6s1_stb),
    .s1_we_o(m6s1_we),
    .s2_ack_i(m6s2_ack),
    .s2_addr_o(m6s2_addr),
    .s2_cyc_o(m6s2_cyc),
    .s2_data_i(m6s2_data_i),
    .s2_data_o(m6s2_data_o),
    .s2_err_i(m6s2_err),
    .s2_rty_i(m6s2_rty),
    .s2_sel_o(m6s2_sel),
    .s2_stb_o(m6s2_stb),
    .s2_we_o(m6s2_we),
    .s3_ack_i(m6s3_ack),
    .s3_addr_o(m6s3_addr),
    .s3_cyc_o(m6s3_cyc),
    .s3_data_i(m6s3_data_i),
    .s3_data_o(m6s3_data_o),
    .s3_err_i(m6s3_err),
    .s3_rty_i(m6s3_rty),
    .s3_sel_o(m6s3_sel),
    .s3_stb_o(m6s3_stb),
    .s3_we_o(m6s3_we),
    .s4_ack_i(m6s4_ack),
    .s4_addr_o(m6s4_addr),
    .s4_cyc_o(m6s4_cyc),
    .s4_data_i(m6s4_data_i),
    .s4_data_o(m6s4_data_o),
    .s4_err_i(m6s4_err),
    .s4_rty_i(m6s4_rty),
    .s4_sel_o(m6s4_sel),
    .s4_stb_o(m6s4_stb),
    .s4_we_o(m6s4_we),
    .s5_ack_i(m6s5_ack),
    .s5_addr_o(m6s5_addr),
    .s5_cyc_o(m6s5_cyc),
    .s5_data_i(m6s5_data_i),
    .s5_data_o(m6s5_data_o),
    .s5_err_i(m6s5_err),
    .s5_rty_i(m6s5_rty),
    .s5_sel_o(m6s5_sel),
    .s5_stb_o(m6s5_stb),
    .s5_we_o(m6s5_we),
    .s6_ack_i(m6s6_ack),
    .s6_addr_o(m6s6_addr),
    .s6_cyc_o(m6s6_cyc),
    .s6_data_i(m6s6_data_i),
    .s6_data_o(m6s6_data_o),
    .s6_err_i(m6s6_err),
    .s6_rty_i(m6s6_rty),
    .s6_sel_o(m6s6_sel),
    .s6_stb_o(m6s6_stb),
    .s6_we_o(m6s6_we),
    .s7_ack_i(m6s7_ack),
    .s7_addr_o(m6s7_addr),
    .s7_cyc_o(m6s7_cyc),
    .s7_data_i(m6s7_data_i),
    .s7_data_o(m6s7_data_o),
    .s7_err_i(m6s7_err),
    .s7_rty_i(m6s7_rty),
    .s7_sel_o(m6s7_sel),
    .s7_stb_o(m6s7_stb),
    .s7_we_o(m6s7_we),
    .s8_ack_i(m6s8_ack),
    .s8_addr_o(m6s8_addr),
    .s8_cyc_o(m6s8_cyc),
    .s8_data_i(m6s8_data_i),
    .s8_data_o(m6s8_data_o),
    .s8_err_i(m6s8_err),
    .s8_rty_i(m6s8_rty),
    .s8_sel_o(m6s8_sel),
    .s8_stb_o(m6s8_stb),
    .s8_we_o(m6s8_we),
    .s9_ack_i(m6s9_ack),
    .s9_addr_o(m6s9_addr),
    .s9_cyc_o(m6s9_cyc),
    .s9_data_i(m6s9_data_i),
    .s9_data_o(m6s9_data_o),
    .s9_err_i(m6s9_err),
    .s9_rty_i(m6s9_rty),
    .s9_sel_o(m6s9_sel),
    .s9_stb_o(m6s9_stb),
    .s9_we_o(m6s9_we),
    .wb_ack_o(_0062_),
    .wb_addr_i(_0063_),
    .wb_cyc_i(_0064_),
    .wb_data_i(_0065_),
    .wb_data_o(_0066_),
    .wb_err_o(_0067_),
    .wb_rty_o(_0068_),
    .wb_sel_i(_0069_),
    .wb_stb_i(_0070_),
    .wb_we_i(_0071_)
  );
\$paramod$7ef9a024e49224e54bf5d1f376214065d47809cb\wb_conmax_master_if   m7 (
    .clk_i(_0001_),
    .rst_i(_0082_),
    .s0_ack_i(m7s0_ack),
    .s0_addr_o(m7s0_addr),
    .s0_cyc_o(m7s0_cyc),
    .s0_data_i(m7s0_data_i),
    .s0_data_o(m7s0_data_o),
    .s0_err_i(m7s0_err),
    .s0_rty_i(m7s0_rty),
    .s0_sel_o(m7s0_sel),
    .s0_stb_o(m7s0_stb),
    .s0_we_o(m7s0_we),
    .s10_ack_i(m7s10_ack),
    .s10_addr_o(m7s10_addr),
    .s10_cyc_o(m7s10_cyc),
    .s10_data_i(m7s10_data_i),
    .s10_data_o(m7s10_data_o),
    .s10_err_i(m7s10_err),
    .s10_rty_i(m7s10_rty),
    .s10_sel_o(m7s10_sel),
    .s10_stb_o(m7s10_stb),
    .s10_we_o(m7s10_we),
    .s11_ack_i(m7s11_ack),
    .s11_addr_o(m7s11_addr),
    .s11_cyc_o(m7s11_cyc),
    .s11_data_i(m7s11_data_i),
    .s11_data_o(m7s11_data_o),
    .s11_err_i(m7s11_err),
    .s11_rty_i(m7s11_rty),
    .s11_sel_o(m7s11_sel),
    .s11_stb_o(m7s11_stb),
    .s11_we_o(m7s11_we),
    .s12_ack_i(m7s12_ack),
    .s12_addr_o(m7s12_addr),
    .s12_cyc_o(m7s12_cyc),
    .s12_data_i(m7s12_data_i),
    .s12_data_o(m7s12_data_o),
    .s12_err_i(m7s12_err),
    .s12_rty_i(m7s12_rty),
    .s12_sel_o(m7s12_sel),
    .s12_stb_o(m7s12_stb),
    .s12_we_o(m7s12_we),
    .s13_ack_i(m7s13_ack),
    .s13_addr_o(m7s13_addr),
    .s13_cyc_o(m7s13_cyc),
    .s13_data_i(m7s13_data_i),
    .s13_data_o(m7s13_data_o),
    .s13_err_i(m7s13_err),
    .s13_rty_i(m7s13_rty),
    .s13_sel_o(m7s13_sel),
    .s13_stb_o(m7s13_stb),
    .s13_we_o(m7s13_we),
    .s14_ack_i(m7s14_ack),
    .s14_addr_o(m7s14_addr),
    .s14_cyc_o(m7s14_cyc),
    .s14_data_i(m7s14_data_i),
    .s14_data_o(m7s14_data_o),
    .s14_err_i(m7s14_err),
    .s14_rty_i(m7s14_rty),
    .s14_sel_o(m7s14_sel),
    .s14_stb_o(m7s14_stb),
    .s14_we_o(m7s14_we),
    .s15_ack_i(m7s15_ack),
    .s15_addr_o(m7s15_addr),
    .s15_cyc_o(m7s15_cyc),
    .s15_data_i(m7s15_data_i),
    .s15_data_o(m7s15_data_o),
    .s15_err_i(m7s15_err),
    .s15_rty_i(m7s15_rty),
    .s15_sel_o(m7s15_sel),
    .s15_stb_o(m7s15_stb),
    .s15_we_o(m7s15_we),
    .s1_ack_i(m7s1_ack),
    .s1_addr_o(m7s1_addr),
    .s1_cyc_o(m7s1_cyc),
    .s1_data_i(m7s1_data_i),
    .s1_data_o(m7s1_data_o),
    .s1_err_i(m7s1_err),
    .s1_rty_i(m7s1_rty),
    .s1_sel_o(m7s1_sel),
    .s1_stb_o(m7s1_stb),
    .s1_we_o(m7s1_we),
    .s2_ack_i(m7s2_ack),
    .s2_addr_o(m7s2_addr),
    .s2_cyc_o(m7s2_cyc),
    .s2_data_i(m7s2_data_i),
    .s2_data_o(m7s2_data_o),
    .s2_err_i(m7s2_err),
    .s2_rty_i(m7s2_rty),
    .s2_sel_o(m7s2_sel),
    .s2_stb_o(m7s2_stb),
    .s2_we_o(m7s2_we),
    .s3_ack_i(m7s3_ack),
    .s3_addr_o(m7s3_addr),
    .s3_cyc_o(m7s3_cyc),
    .s3_data_i(m7s3_data_i),
    .s3_data_o(m7s3_data_o),
    .s3_err_i(m7s3_err),
    .s3_rty_i(m7s3_rty),
    .s3_sel_o(m7s3_sel),
    .s3_stb_o(m7s3_stb),
    .s3_we_o(m7s3_we),
    .s4_ack_i(m7s4_ack),
    .s4_addr_o(m7s4_addr),
    .s4_cyc_o(m7s4_cyc),
    .s4_data_i(m7s4_data_i),
    .s4_data_o(m7s4_data_o),
    .s4_err_i(m7s4_err),
    .s4_rty_i(m7s4_rty),
    .s4_sel_o(m7s4_sel),
    .s4_stb_o(m7s4_stb),
    .s4_we_o(m7s4_we),
    .s5_ack_i(m7s5_ack),
    .s5_addr_o(m7s5_addr),
    .s5_cyc_o(m7s5_cyc),
    .s5_data_i(m7s5_data_i),
    .s5_data_o(m7s5_data_o),
    .s5_err_i(m7s5_err),
    .s5_rty_i(m7s5_rty),
    .s5_sel_o(m7s5_sel),
    .s5_stb_o(m7s5_stb),
    .s5_we_o(m7s5_we),
    .s6_ack_i(m7s6_ack),
    .s6_addr_o(m7s6_addr),
    .s6_cyc_o(m7s6_cyc),
    .s6_data_i(m7s6_data_i),
    .s6_data_o(m7s6_data_o),
    .s6_err_i(m7s6_err),
    .s6_rty_i(m7s6_rty),
    .s6_sel_o(m7s6_sel),
    .s6_stb_o(m7s6_stb),
    .s6_we_o(m7s6_we),
    .s7_ack_i(m7s7_ack),
    .s7_addr_o(m7s7_addr),
    .s7_cyc_o(m7s7_cyc),
    .s7_data_i(m7s7_data_i),
    .s7_data_o(m7s7_data_o),
    .s7_err_i(m7s7_err),
    .s7_rty_i(m7s7_rty),
    .s7_sel_o(m7s7_sel),
    .s7_stb_o(m7s7_stb),
    .s7_we_o(m7s7_we),
    .s8_ack_i(m7s8_ack),
    .s8_addr_o(m7s8_addr),
    .s8_cyc_o(m7s8_cyc),
    .s8_data_i(m7s8_data_i),
    .s8_data_o(m7s8_data_o),
    .s8_err_i(m7s8_err),
    .s8_rty_i(m7s8_rty),
    .s8_sel_o(m7s8_sel),
    .s8_stb_o(m7s8_stb),
    .s8_we_o(m7s8_we),
    .s9_ack_i(m7s9_ack),
    .s9_addr_o(m7s9_addr),
    .s9_cyc_o(m7s9_cyc),
    .s9_data_i(m7s9_data_i),
    .s9_data_o(m7s9_data_o),
    .s9_err_i(m7s9_err),
    .s9_rty_i(m7s9_rty),
    .s9_sel_o(m7s9_sel),
    .s9_stb_o(m7s9_stb),
    .s9_we_o(m7s9_we),
    .wb_ack_o(_0072_),
    .wb_addr_i(_0073_),
    .wb_cyc_i(_0074_),
    .wb_data_i(_0075_),
    .wb_data_o(_0076_),
    .wb_err_o(_0077_),
    .wb_rty_o(_0078_),
    .wb_sel_i(_0079_),
    .wb_stb_i(_0080_),
    .wb_we_i(_0081_)
  );
\$paramod$9dc2a30a66a5cd1c6354168b9c37f048ec339685\wb_conmax_rf   rf (
    .clk_i(_0001_),
    .conf0(conf0),
    .conf1(conf1),
    .conf10(conf10),
    .conf11(conf11),
    .conf12(conf12),
    .conf13(conf13),
    .conf14(conf14),
    .conf15(conf15),
    .conf2(conf2),
    .conf3(conf3),
    .conf4(conf4),
    .conf5(conf5),
    .conf6(conf6),
    .conf7(conf7),
    .conf8(conf8),
    .conf9(conf9),
    .e_wb_ack_i(_0143_),
    .e_wb_addr_o(_0144_),
    .e_wb_cyc_o(_0145_),
    .e_wb_data_i(_0146_),
    .e_wb_data_o(_0147_),
    .e_wb_err_i(_0148_),
    .e_wb_rty_i(_0149_),
    .e_wb_sel_o(_0150_),
    .e_wb_stb_o(_0151_),
    .e_wb_we_o(_0152_),
    .i_wb_ack_o(i_s15_ack_i),
    .i_wb_addr_i(i_s15_addr_o),
    .i_wb_cyc_i(i_s15_cyc_o),
    .i_wb_data_i(i_s15_data_o),
    .i_wb_data_o(i_s15_data_i),
    .i_wb_err_o(i_s15_err_i),
    .i_wb_rty_o(i_s15_rty_i),
    .i_wb_sel_i(i_s15_sel_o),
    .i_wb_stb_i(i_s15_stb_o),
    .i_wb_we_i(i_s15_we_o),
    .rst_i(_0082_)
  );
\$paramod$babc7f28591f52523637895ab98a5c04b5a93873\wb_conmax_slave_if   s0 (
    .clk_i(_0001_),
    .conf(conf0),
    .m0_ack_o(m0s0_ack),
    .m0_addr_i(m0s0_addr),
    .m0_cyc_i(m0s0_cyc),
    .m0_data_i(m0s0_data_o),
    .m0_data_o(m0s0_data_i),
    .m0_err_o(m0s0_err),
    .m0_rty_o(m0s0_rty),
    .m0_sel_i(m0s0_sel),
    .m0_stb_i(m0s0_stb),
    .m0_we_i(m0s0_we),
    .m1_ack_o(m1s0_ack),
    .m1_addr_i(m1s0_addr),
    .m1_cyc_i(m1s0_cyc),
    .m1_data_i(m1s0_data_o),
    .m1_data_o(m1s0_data_i),
    .m1_err_o(m1s0_err),
    .m1_rty_o(m1s0_rty),
    .m1_sel_i(m1s0_sel),
    .m1_stb_i(m1s0_stb),
    .m1_we_i(m1s0_we),
    .m2_ack_o(m2s0_ack),
    .m2_addr_i(m2s0_addr),
    .m2_cyc_i(m2s0_cyc),
    .m2_data_i(m2s0_data_o),
    .m2_data_o(m2s0_data_i),
    .m2_err_o(m2s0_err),
    .m2_rty_o(m2s0_rty),
    .m2_sel_i(m2s0_sel),
    .m2_stb_i(m2s0_stb),
    .m2_we_i(m2s0_we),
    .m3_ack_o(m3s0_ack),
    .m3_addr_i(m3s0_addr),
    .m3_cyc_i(m3s0_cyc),
    .m3_data_i(m3s0_data_o),
    .m3_data_o(m3s0_data_i),
    .m3_err_o(m3s0_err),
    .m3_rty_o(m3s0_rty),
    .m3_sel_i(m3s0_sel),
    .m3_stb_i(m3s0_stb),
    .m3_we_i(m3s0_we),
    .m4_ack_o(m4s0_ack),
    .m4_addr_i(m4s0_addr),
    .m4_cyc_i(m4s0_cyc),
    .m4_data_i(m4s0_data_o),
    .m4_data_o(m4s0_data_i),
    .m4_err_o(m4s0_err),
    .m4_rty_o(m4s0_rty),
    .m4_sel_i(m4s0_sel),
    .m4_stb_i(m4s0_stb),
    .m4_we_i(m4s0_we),
    .m5_ack_o(m5s0_ack),
    .m5_addr_i(m5s0_addr),
    .m5_cyc_i(m5s0_cyc),
    .m5_data_i(m5s0_data_o),
    .m5_data_o(m5s0_data_i),
    .m5_err_o(m5s0_err),
    .m5_rty_o(m5s0_rty),
    .m5_sel_i(m5s0_sel),
    .m5_stb_i(m5s0_stb),
    .m5_we_i(m5s0_we),
    .m6_ack_o(m6s0_ack),
    .m6_addr_i(m6s0_addr),
    .m6_cyc_i(m6s0_cyc),
    .m6_data_i(m6s0_data_o),
    .m6_data_o(m6s0_data_i),
    .m6_err_o(m6s0_err),
    .m6_rty_o(m6s0_rty),
    .m6_sel_i(m6s0_sel),
    .m6_stb_i(m6s0_stb),
    .m6_we_i(m6s0_we),
    .m7_ack_o(m7s0_ack),
    .m7_addr_i(m7s0_addr),
    .m7_cyc_i(m7s0_cyc),
    .m7_data_i(m7s0_data_o),
    .m7_data_o(m7s0_data_i),
    .m7_err_o(m7s0_err),
    .m7_rty_o(m7s0_rty),
    .m7_sel_i(m7s0_sel),
    .m7_stb_i(m7s0_stb),
    .m7_we_i(m7s0_we),
    .rst_i(_0082_),
    .wb_ack_i(_0083_),
    .wb_addr_o(_0084_),
    .wb_cyc_o(_0085_),
    .wb_data_i(_0086_),
    .wb_data_o(_0087_),
    .wb_err_i(_0088_),
    .wb_rty_i(_0089_),
    .wb_sel_o(_0090_),
    .wb_stb_o(_0091_),
    .wb_we_o(_0092_)
  );
\$paramod$babc7f28591f52523637895ab98a5c04b5a93873\wb_conmax_slave_if   s1 (
    .clk_i(_0001_),
    .conf(conf1),
    .m0_ack_o(m0s1_ack),
    .m0_addr_i(m0s1_addr),
    .m0_cyc_i(m0s1_cyc),
    .m0_data_i(m0s1_data_o),
    .m0_data_o(m0s1_data_i),
    .m0_err_o(m0s1_err),
    .m0_rty_o(m0s1_rty),
    .m0_sel_i(m0s1_sel),
    .m0_stb_i(m0s1_stb),
    .m0_we_i(m0s1_we),
    .m1_ack_o(m1s1_ack),
    .m1_addr_i(m1s1_addr),
    .m1_cyc_i(m1s1_cyc),
    .m1_data_i(m1s1_data_o),
    .m1_data_o(m1s1_data_i),
    .m1_err_o(m1s1_err),
    .m1_rty_o(m1s1_rty),
    .m1_sel_i(m1s1_sel),
    .m1_stb_i(m1s1_stb),
    .m1_we_i(m1s1_we),
    .m2_ack_o(m2s1_ack),
    .m2_addr_i(m2s1_addr),
    .m2_cyc_i(m2s1_cyc),
    .m2_data_i(m2s1_data_o),
    .m2_data_o(m2s1_data_i),
    .m2_err_o(m2s1_err),
    .m2_rty_o(m2s1_rty),
    .m2_sel_i(m2s1_sel),
    .m2_stb_i(m2s1_stb),
    .m2_we_i(m2s1_we),
    .m3_ack_o(m3s1_ack),
    .m3_addr_i(m3s1_addr),
    .m3_cyc_i(m3s1_cyc),
    .m3_data_i(m3s1_data_o),
    .m3_data_o(m3s1_data_i),
    .m3_err_o(m3s1_err),
    .m3_rty_o(m3s1_rty),
    .m3_sel_i(m3s1_sel),
    .m3_stb_i(m3s1_stb),
    .m3_we_i(m3s1_we),
    .m4_ack_o(m4s1_ack),
    .m4_addr_i(m4s1_addr),
    .m4_cyc_i(m4s1_cyc),
    .m4_data_i(m4s1_data_o),
    .m4_data_o(m4s1_data_i),
    .m4_err_o(m4s1_err),
    .m4_rty_o(m4s1_rty),
    .m4_sel_i(m4s1_sel),
    .m4_stb_i(m4s1_stb),
    .m4_we_i(m4s1_we),
    .m5_ack_o(m5s1_ack),
    .m5_addr_i(m5s1_addr),
    .m5_cyc_i(m5s1_cyc),
    .m5_data_i(m5s1_data_o),
    .m5_data_o(m5s1_data_i),
    .m5_err_o(m5s1_err),
    .m5_rty_o(m5s1_rty),
    .m5_sel_i(m5s1_sel),
    .m5_stb_i(m5s1_stb),
    .m5_we_i(m5s1_we),
    .m6_ack_o(m6s1_ack),
    .m6_addr_i(m6s1_addr),
    .m6_cyc_i(m6s1_cyc),
    .m6_data_i(m6s1_data_o),
    .m6_data_o(m6s1_data_i),
    .m6_err_o(m6s1_err),
    .m6_rty_o(m6s1_rty),
    .m6_sel_i(m6s1_sel),
    .m6_stb_i(m6s1_stb),
    .m6_we_i(m6s1_we),
    .m7_ack_o(m7s1_ack),
    .m7_addr_i(m7s1_addr),
    .m7_cyc_i(m7s1_cyc),
    .m7_data_i(m7s1_data_o),
    .m7_data_o(m7s1_data_i),
    .m7_err_o(m7s1_err),
    .m7_rty_o(m7s1_rty),
    .m7_sel_i(m7s1_sel),
    .m7_stb_i(m7s1_stb),
    .m7_we_i(m7s1_we),
    .rst_i(_0082_),
    .wb_ack_i(_0153_),
    .wb_addr_o(_0154_),
    .wb_cyc_o(_0155_),
    .wb_data_i(_0156_),
    .wb_data_o(_0157_),
    .wb_err_i(_0158_),
    .wb_rty_i(_0159_),
    .wb_sel_o(_0160_),
    .wb_stb_o(_0161_),
    .wb_we_o(_0162_)
  );
\$paramod$babc7f28591f52523637895ab98a5c04b5a93873\wb_conmax_slave_if   s10 (
    .clk_i(_0001_),
    .conf(conf10),
    .m0_ack_o(m0s10_ack),
    .m0_addr_i(m0s10_addr),
    .m0_cyc_i(m0s10_cyc),
    .m0_data_i(m0s10_data_o),
    .m0_data_o(m0s10_data_i),
    .m0_err_o(m0s10_err),
    .m0_rty_o(m0s10_rty),
    .m0_sel_i(m0s10_sel),
    .m0_stb_i(m0s10_stb),
    .m0_we_i(m0s10_we),
    .m1_ack_o(m1s10_ack),
    .m1_addr_i(m1s10_addr),
    .m1_cyc_i(m1s10_cyc),
    .m1_data_i(m1s10_data_o),
    .m1_data_o(m1s10_data_i),
    .m1_err_o(m1s10_err),
    .m1_rty_o(m1s10_rty),
    .m1_sel_i(m1s10_sel),
    .m1_stb_i(m1s10_stb),
    .m1_we_i(m1s10_we),
    .m2_ack_o(m2s10_ack),
    .m2_addr_i(m2s10_addr),
    .m2_cyc_i(m2s10_cyc),
    .m2_data_i(m2s10_data_o),
    .m2_data_o(m2s10_data_i),
    .m2_err_o(m2s10_err),
    .m2_rty_o(m2s10_rty),
    .m2_sel_i(m2s10_sel),
    .m2_stb_i(m2s10_stb),
    .m2_we_i(m2s10_we),
    .m3_ack_o(m3s10_ack),
    .m3_addr_i(m3s10_addr),
    .m3_cyc_i(m3s10_cyc),
    .m3_data_i(m3s10_data_o),
    .m3_data_o(m3s10_data_i),
    .m3_err_o(m3s10_err),
    .m3_rty_o(m3s10_rty),
    .m3_sel_i(m3s10_sel),
    .m3_stb_i(m3s10_stb),
    .m3_we_i(m3s10_we),
    .m4_ack_o(m4s10_ack),
    .m4_addr_i(m4s10_addr),
    .m4_cyc_i(m4s10_cyc),
    .m4_data_i(m4s10_data_o),
    .m4_data_o(m4s10_data_i),
    .m4_err_o(m4s10_err),
    .m4_rty_o(m4s10_rty),
    .m4_sel_i(m4s10_sel),
    .m4_stb_i(m4s10_stb),
    .m4_we_i(m4s10_we),
    .m5_ack_o(m5s10_ack),
    .m5_addr_i(m5s10_addr),
    .m5_cyc_i(m5s10_cyc),
    .m5_data_i(m5s10_data_o),
    .m5_data_o(m5s10_data_i),
    .m5_err_o(m5s10_err),
    .m5_rty_o(m5s10_rty),
    .m5_sel_i(m5s10_sel),
    .m5_stb_i(m5s10_stb),
    .m5_we_i(m5s10_we),
    .m6_ack_o(m6s10_ack),
    .m6_addr_i(m6s10_addr),
    .m6_cyc_i(m6s10_cyc),
    .m6_data_i(m6s10_data_o),
    .m6_data_o(m6s10_data_i),
    .m6_err_o(m6s10_err),
    .m6_rty_o(m6s10_rty),
    .m6_sel_i(m6s10_sel),
    .m6_stb_i(m6s10_stb),
    .m6_we_i(m6s10_we),
    .m7_ack_o(m7s10_ack),
    .m7_addr_i(m7s10_addr),
    .m7_cyc_i(m7s10_cyc),
    .m7_data_i(m7s10_data_o),
    .m7_data_o(m7s10_data_i),
    .m7_err_o(m7s10_err),
    .m7_rty_o(m7s10_rty),
    .m7_sel_i(m7s10_sel),
    .m7_stb_i(m7s10_stb),
    .m7_we_i(m7s10_we),
    .rst_i(_0082_),
    .wb_ack_i(_0093_),
    .wb_addr_o(_0094_),
    .wb_cyc_o(_0095_),
    .wb_data_i(_0096_),
    .wb_data_o(_0097_),
    .wb_err_i(_0098_),
    .wb_rty_i(_0099_),
    .wb_sel_o(_0100_),
    .wb_stb_o(_0101_),
    .wb_we_o(_0102_)
  );
\$paramod$babc7f28591f52523637895ab98a5c04b5a93873\wb_conmax_slave_if   s11 (
    .clk_i(_0001_),
    .conf(conf11),
    .m0_ack_o(m0s11_ack),
    .m0_addr_i(m0s11_addr),
    .m0_cyc_i(m0s11_cyc),
    .m0_data_i(m0s11_data_o),
    .m0_data_o(m0s11_data_i),
    .m0_err_o(m0s11_err),
    .m0_rty_o(m0s11_rty),
    .m0_sel_i(m0s11_sel),
    .m0_stb_i(m0s11_stb),
    .m0_we_i(m0s11_we),
    .m1_ack_o(m1s11_ack),
    .m1_addr_i(m1s11_addr),
    .m1_cyc_i(m1s11_cyc),
    .m1_data_i(m1s11_data_o),
    .m1_data_o(m1s11_data_i),
    .m1_err_o(m1s11_err),
    .m1_rty_o(m1s11_rty),
    .m1_sel_i(m1s11_sel),
    .m1_stb_i(m1s11_stb),
    .m1_we_i(m1s11_we),
    .m2_ack_o(m2s11_ack),
    .m2_addr_i(m2s11_addr),
    .m2_cyc_i(m2s11_cyc),
    .m2_data_i(m2s11_data_o),
    .m2_data_o(m2s11_data_i),
    .m2_err_o(m2s11_err),
    .m2_rty_o(m2s11_rty),
    .m2_sel_i(m2s11_sel),
    .m2_stb_i(m2s11_stb),
    .m2_we_i(m2s11_we),
    .m3_ack_o(m3s11_ack),
    .m3_addr_i(m3s11_addr),
    .m3_cyc_i(m3s11_cyc),
    .m3_data_i(m3s11_data_o),
    .m3_data_o(m3s11_data_i),
    .m3_err_o(m3s11_err),
    .m3_rty_o(m3s11_rty),
    .m3_sel_i(m3s11_sel),
    .m3_stb_i(m3s11_stb),
    .m3_we_i(m3s11_we),
    .m4_ack_o(m4s11_ack),
    .m4_addr_i(m4s11_addr),
    .m4_cyc_i(m4s11_cyc),
    .m4_data_i(m4s11_data_o),
    .m4_data_o(m4s11_data_i),
    .m4_err_o(m4s11_err),
    .m4_rty_o(m4s11_rty),
    .m4_sel_i(m4s11_sel),
    .m4_stb_i(m4s11_stb),
    .m4_we_i(m4s11_we),
    .m5_ack_o(m5s11_ack),
    .m5_addr_i(m5s11_addr),
    .m5_cyc_i(m5s11_cyc),
    .m5_data_i(m5s11_data_o),
    .m5_data_o(m5s11_data_i),
    .m5_err_o(m5s11_err),
    .m5_rty_o(m5s11_rty),
    .m5_sel_i(m5s11_sel),
    .m5_stb_i(m5s11_stb),
    .m5_we_i(m5s11_we),
    .m6_ack_o(m6s11_ack),
    .m6_addr_i(m6s11_addr),
    .m6_cyc_i(m6s11_cyc),
    .m6_data_i(m6s11_data_o),
    .m6_data_o(m6s11_data_i),
    .m6_err_o(m6s11_err),
    .m6_rty_o(m6s11_rty),
    .m6_sel_i(m6s11_sel),
    .m6_stb_i(m6s11_stb),
    .m6_we_i(m6s11_we),
    .m7_ack_o(m7s11_ack),
    .m7_addr_i(m7s11_addr),
    .m7_cyc_i(m7s11_cyc),
    .m7_data_i(m7s11_data_o),
    .m7_data_o(m7s11_data_i),
    .m7_err_o(m7s11_err),
    .m7_rty_o(m7s11_rty),
    .m7_sel_i(m7s11_sel),
    .m7_stb_i(m7s11_stb),
    .m7_we_i(m7s11_we),
    .rst_i(_0082_),
    .wb_ack_i(_0103_),
    .wb_addr_o(_0104_),
    .wb_cyc_o(_0105_),
    .wb_data_i(_0106_),
    .wb_data_o(_0107_),
    .wb_err_i(_0108_),
    .wb_rty_i(_0109_),
    .wb_sel_o(_0110_),
    .wb_stb_o(_0111_),
    .wb_we_o(_0112_)
  );
\$paramod$babc7f28591f52523637895ab98a5c04b5a93873\wb_conmax_slave_if   s12 (
    .clk_i(_0001_),
    .conf(conf12),
    .m0_ack_o(m0s12_ack),
    .m0_addr_i(m0s12_addr),
    .m0_cyc_i(m0s12_cyc),
    .m0_data_i(m0s12_data_o),
    .m0_data_o(m0s12_data_i),
    .m0_err_o(m0s12_err),
    .m0_rty_o(m0s12_rty),
    .m0_sel_i(m0s12_sel),
    .m0_stb_i(m0s12_stb),
    .m0_we_i(m0s12_we),
    .m1_ack_o(m1s12_ack),
    .m1_addr_i(m1s12_addr),
    .m1_cyc_i(m1s12_cyc),
    .m1_data_i(m1s12_data_o),
    .m1_data_o(m1s12_data_i),
    .m1_err_o(m1s12_err),
    .m1_rty_o(m1s12_rty),
    .m1_sel_i(m1s12_sel),
    .m1_stb_i(m1s12_stb),
    .m1_we_i(m1s12_we),
    .m2_ack_o(m2s12_ack),
    .m2_addr_i(m2s12_addr),
    .m2_cyc_i(m2s12_cyc),
    .m2_data_i(m2s12_data_o),
    .m2_data_o(m2s12_data_i),
    .m2_err_o(m2s12_err),
    .m2_rty_o(m2s12_rty),
    .m2_sel_i(m2s12_sel),
    .m2_stb_i(m2s12_stb),
    .m2_we_i(m2s12_we),
    .m3_ack_o(m3s12_ack),
    .m3_addr_i(m3s12_addr),
    .m3_cyc_i(m3s12_cyc),
    .m3_data_i(m3s12_data_o),
    .m3_data_o(m3s12_data_i),
    .m3_err_o(m3s12_err),
    .m3_rty_o(m3s12_rty),
    .m3_sel_i(m3s12_sel),
    .m3_stb_i(m3s12_stb),
    .m3_we_i(m3s12_we),
    .m4_ack_o(m4s12_ack),
    .m4_addr_i(m4s12_addr),
    .m4_cyc_i(m4s12_cyc),
    .m4_data_i(m4s12_data_o),
    .m4_data_o(m4s12_data_i),
    .m4_err_o(m4s12_err),
    .m4_rty_o(m4s12_rty),
    .m4_sel_i(m4s12_sel),
    .m4_stb_i(m4s12_stb),
    .m4_we_i(m4s12_we),
    .m5_ack_o(m5s12_ack),
    .m5_addr_i(m5s12_addr),
    .m5_cyc_i(m5s12_cyc),
    .m5_data_i(m5s12_data_o),
    .m5_data_o(m5s12_data_i),
    .m5_err_o(m5s12_err),
    .m5_rty_o(m5s12_rty),
    .m5_sel_i(m5s12_sel),
    .m5_stb_i(m5s12_stb),
    .m5_we_i(m5s12_we),
    .m6_ack_o(m6s12_ack),
    .m6_addr_i(m6s12_addr),
    .m6_cyc_i(m6s12_cyc),
    .m6_data_i(m6s12_data_o),
    .m6_data_o(m6s12_data_i),
    .m6_err_o(m6s12_err),
    .m6_rty_o(m6s12_rty),
    .m6_sel_i(m6s12_sel),
    .m6_stb_i(m6s12_stb),
    .m6_we_i(m6s12_we),
    .m7_ack_o(m7s12_ack),
    .m7_addr_i(m7s12_addr),
    .m7_cyc_i(m7s12_cyc),
    .m7_data_i(m7s12_data_o),
    .m7_data_o(m7s12_data_i),
    .m7_err_o(m7s12_err),
    .m7_rty_o(m7s12_rty),
    .m7_sel_i(m7s12_sel),
    .m7_stb_i(m7s12_stb),
    .m7_we_i(m7s12_we),
    .rst_i(_0082_),
    .wb_ack_i(_0113_),
    .wb_addr_o(_0114_),
    .wb_cyc_o(_0115_),
    .wb_data_i(_0116_),
    .wb_data_o(_0117_),
    .wb_err_i(_0118_),
    .wb_rty_i(_0119_),
    .wb_sel_o(_0120_),
    .wb_stb_o(_0121_),
    .wb_we_o(_0122_)
  );
\$paramod$babc7f28591f52523637895ab98a5c04b5a93873\wb_conmax_slave_if   s13 (
    .clk_i(_0001_),
    .conf(conf13),
    .m0_ack_o(m0s13_ack),
    .m0_addr_i(m0s13_addr),
    .m0_cyc_i(m0s13_cyc),
    .m0_data_i(m0s13_data_o),
    .m0_data_o(m0s13_data_i),
    .m0_err_o(m0s13_err),
    .m0_rty_o(m0s13_rty),
    .m0_sel_i(m0s13_sel),
    .m0_stb_i(m0s13_stb),
    .m0_we_i(m0s13_we),
    .m1_ack_o(m1s13_ack),
    .m1_addr_i(m1s13_addr),
    .m1_cyc_i(m1s13_cyc),
    .m1_data_i(m1s13_data_o),
    .m1_data_o(m1s13_data_i),
    .m1_err_o(m1s13_err),
    .m1_rty_o(m1s13_rty),
    .m1_sel_i(m1s13_sel),
    .m1_stb_i(m1s13_stb),
    .m1_we_i(m1s13_we),
    .m2_ack_o(m2s13_ack),
    .m2_addr_i(m2s13_addr),
    .m2_cyc_i(m2s13_cyc),
    .m2_data_i(m2s13_data_o),
    .m2_data_o(m2s13_data_i),
    .m2_err_o(m2s13_err),
    .m2_rty_o(m2s13_rty),
    .m2_sel_i(m2s13_sel),
    .m2_stb_i(m2s13_stb),
    .m2_we_i(m2s13_we),
    .m3_ack_o(m3s13_ack),
    .m3_addr_i(m3s13_addr),
    .m3_cyc_i(m3s13_cyc),
    .m3_data_i(m3s13_data_o),
    .m3_data_o(m3s13_data_i),
    .m3_err_o(m3s13_err),
    .m3_rty_o(m3s13_rty),
    .m3_sel_i(m3s13_sel),
    .m3_stb_i(m3s13_stb),
    .m3_we_i(m3s13_we),
    .m4_ack_o(m4s13_ack),
    .m4_addr_i(m4s13_addr),
    .m4_cyc_i(m4s13_cyc),
    .m4_data_i(m4s13_data_o),
    .m4_data_o(m4s13_data_i),
    .m4_err_o(m4s13_err),
    .m4_rty_o(m4s13_rty),
    .m4_sel_i(m4s13_sel),
    .m4_stb_i(m4s13_stb),
    .m4_we_i(m4s13_we),
    .m5_ack_o(m5s13_ack),
    .m5_addr_i(m5s13_addr),
    .m5_cyc_i(m5s13_cyc),
    .m5_data_i(m5s13_data_o),
    .m5_data_o(m5s13_data_i),
    .m5_err_o(m5s13_err),
    .m5_rty_o(m5s13_rty),
    .m5_sel_i(m5s13_sel),
    .m5_stb_i(m5s13_stb),
    .m5_we_i(m5s13_we),
    .m6_ack_o(m6s13_ack),
    .m6_addr_i(m6s13_addr),
    .m6_cyc_i(m6s13_cyc),
    .m6_data_i(m6s13_data_o),
    .m6_data_o(m6s13_data_i),
    .m6_err_o(m6s13_err),
    .m6_rty_o(m6s13_rty),
    .m6_sel_i(m6s13_sel),
    .m6_stb_i(m6s13_stb),
    .m6_we_i(m6s13_we),
    .m7_ack_o(m7s13_ack),
    .m7_addr_i(m7s13_addr),
    .m7_cyc_i(m7s13_cyc),
    .m7_data_i(m7s13_data_o),
    .m7_data_o(m7s13_data_i),
    .m7_err_o(m7s13_err),
    .m7_rty_o(m7s13_rty),
    .m7_sel_i(m7s13_sel),
    .m7_stb_i(m7s13_stb),
    .m7_we_i(m7s13_we),
    .rst_i(_0082_),
    .wb_ack_i(_0123_),
    .wb_addr_o(_0124_),
    .wb_cyc_o(_0125_),
    .wb_data_i(_0126_),
    .wb_data_o(_0127_),
    .wb_err_i(_0128_),
    .wb_rty_i(_0129_),
    .wb_sel_o(_0130_),
    .wb_stb_o(_0131_),
    .wb_we_o(_0132_)
  );
\$paramod$babc7f28591f52523637895ab98a5c04b5a93873\wb_conmax_slave_if   s14 (
    .clk_i(_0001_),
    .conf(conf14),
    .m0_ack_o(m0s14_ack),
    .m0_addr_i(m0s14_addr),
    .m0_cyc_i(m0s14_cyc),
    .m0_data_i(m0s14_data_o),
    .m0_data_o(m0s14_data_i),
    .m0_err_o(m0s14_err),
    .m0_rty_o(m0s14_rty),
    .m0_sel_i(m0s14_sel),
    .m0_stb_i(m0s14_stb),
    .m0_we_i(m0s14_we),
    .m1_ack_o(m1s14_ack),
    .m1_addr_i(m1s14_addr),
    .m1_cyc_i(m1s14_cyc),
    .m1_data_i(m1s14_data_o),
    .m1_data_o(m1s14_data_i),
    .m1_err_o(m1s14_err),
    .m1_rty_o(m1s14_rty),
    .m1_sel_i(m1s14_sel),
    .m1_stb_i(m1s14_stb),
    .m1_we_i(m1s14_we),
    .m2_ack_o(m2s14_ack),
    .m2_addr_i(m2s14_addr),
    .m2_cyc_i(m2s14_cyc),
    .m2_data_i(m2s14_data_o),
    .m2_data_o(m2s14_data_i),
    .m2_err_o(m2s14_err),
    .m2_rty_o(m2s14_rty),
    .m2_sel_i(m2s14_sel),
    .m2_stb_i(m2s14_stb),
    .m2_we_i(m2s14_we),
    .m3_ack_o(m3s14_ack),
    .m3_addr_i(m3s14_addr),
    .m3_cyc_i(m3s14_cyc),
    .m3_data_i(m3s14_data_o),
    .m3_data_o(m3s14_data_i),
    .m3_err_o(m3s14_err),
    .m3_rty_o(m3s14_rty),
    .m3_sel_i(m3s14_sel),
    .m3_stb_i(m3s14_stb),
    .m3_we_i(m3s14_we),
    .m4_ack_o(m4s14_ack),
    .m4_addr_i(m4s14_addr),
    .m4_cyc_i(m4s14_cyc),
    .m4_data_i(m4s14_data_o),
    .m4_data_o(m4s14_data_i),
    .m4_err_o(m4s14_err),
    .m4_rty_o(m4s14_rty),
    .m4_sel_i(m4s14_sel),
    .m4_stb_i(m4s14_stb),
    .m4_we_i(m4s14_we),
    .m5_ack_o(m5s14_ack),
    .m5_addr_i(m5s14_addr),
    .m5_cyc_i(m5s14_cyc),
    .m5_data_i(m5s14_data_o),
    .m5_data_o(m5s14_data_i),
    .m5_err_o(m5s14_err),
    .m5_rty_o(m5s14_rty),
    .m5_sel_i(m5s14_sel),
    .m5_stb_i(m5s14_stb),
    .m5_we_i(m5s14_we),
    .m6_ack_o(m6s14_ack),
    .m6_addr_i(m6s14_addr),
    .m6_cyc_i(m6s14_cyc),
    .m6_data_i(m6s14_data_o),
    .m6_data_o(m6s14_data_i),
    .m6_err_o(m6s14_err),
    .m6_rty_o(m6s14_rty),
    .m6_sel_i(m6s14_sel),
    .m6_stb_i(m6s14_stb),
    .m6_we_i(m6s14_we),
    .m7_ack_o(m7s14_ack),
    .m7_addr_i(m7s14_addr),
    .m7_cyc_i(m7s14_cyc),
    .m7_data_i(m7s14_data_o),
    .m7_data_o(m7s14_data_i),
    .m7_err_o(m7s14_err),
    .m7_rty_o(m7s14_rty),
    .m7_sel_i(m7s14_sel),
    .m7_stb_i(m7s14_stb),
    .m7_we_i(m7s14_we),
    .rst_i(_0082_),
    .wb_ack_i(_0133_),
    .wb_addr_o(_0134_),
    .wb_cyc_o(_0135_),
    .wb_data_i(_0136_),
    .wb_data_o(_0137_),
    .wb_err_i(_0138_),
    .wb_rty_i(_0139_),
    .wb_sel_o(_0140_),
    .wb_stb_o(_0141_),
    .wb_we_o(_0142_)
  );
\$paramod$babc7f28591f52523637895ab98a5c04b5a93873\wb_conmax_slave_if   s15 (
    .clk_i(_0001_),
    .conf(conf15),
    .m0_ack_o(m0s15_ack),
    .m0_addr_i(m0s15_addr),
    .m0_cyc_i(m0s15_cyc),
    .m0_data_i(m0s15_data_o),
    .m0_data_o(m0s15_data_i),
    .m0_err_o(m0s15_err),
    .m0_rty_o(m0s15_rty),
    .m0_sel_i(m0s15_sel),
    .m0_stb_i(m0s15_stb),
    .m0_we_i(m0s15_we),
    .m1_ack_o(m1s15_ack),
    .m1_addr_i(m1s15_addr),
    .m1_cyc_i(m1s15_cyc),
    .m1_data_i(m1s15_data_o),
    .m1_data_o(m1s15_data_i),
    .m1_err_o(m1s15_err),
    .m1_rty_o(m1s15_rty),
    .m1_sel_i(m1s15_sel),
    .m1_stb_i(m1s15_stb),
    .m1_we_i(m1s15_we),
    .m2_ack_o(m2s15_ack),
    .m2_addr_i(m2s15_addr),
    .m2_cyc_i(m2s15_cyc),
    .m2_data_i(m2s15_data_o),
    .m2_data_o(m2s15_data_i),
    .m2_err_o(m2s15_err),
    .m2_rty_o(m2s15_rty),
    .m2_sel_i(m2s15_sel),
    .m2_stb_i(m2s15_stb),
    .m2_we_i(m2s15_we),
    .m3_ack_o(m3s15_ack),
    .m3_addr_i(m3s15_addr),
    .m3_cyc_i(m3s15_cyc),
    .m3_data_i(m3s15_data_o),
    .m3_data_o(m3s15_data_i),
    .m3_err_o(m3s15_err),
    .m3_rty_o(m3s15_rty),
    .m3_sel_i(m3s15_sel),
    .m3_stb_i(m3s15_stb),
    .m3_we_i(m3s15_we),
    .m4_ack_o(m4s15_ack),
    .m4_addr_i(m4s15_addr),
    .m4_cyc_i(m4s15_cyc),
    .m4_data_i(m4s15_data_o),
    .m4_data_o(m4s15_data_i),
    .m4_err_o(m4s15_err),
    .m4_rty_o(m4s15_rty),
    .m4_sel_i(m4s15_sel),
    .m4_stb_i(m4s15_stb),
    .m4_we_i(m4s15_we),
    .m5_ack_o(m5s15_ack),
    .m5_addr_i(m5s15_addr),
    .m5_cyc_i(m5s15_cyc),
    .m5_data_i(m5s15_data_o),
    .m5_data_o(m5s15_data_i),
    .m5_err_o(m5s15_err),
    .m5_rty_o(m5s15_rty),
    .m5_sel_i(m5s15_sel),
    .m5_stb_i(m5s15_stb),
    .m5_we_i(m5s15_we),
    .m6_ack_o(m6s15_ack),
    .m6_addr_i(m6s15_addr),
    .m6_cyc_i(m6s15_cyc),
    .m6_data_i(m6s15_data_o),
    .m6_data_o(m6s15_data_i),
    .m6_err_o(m6s15_err),
    .m6_rty_o(m6s15_rty),
    .m6_sel_i(m6s15_sel),
    .m6_stb_i(m6s15_stb),
    .m6_we_i(m6s15_we),
    .m7_ack_o(m7s15_ack),
    .m7_addr_i(m7s15_addr),
    .m7_cyc_i(m7s15_cyc),
    .m7_data_i(m7s15_data_o),
    .m7_data_o(m7s15_data_i),
    .m7_err_o(m7s15_err),
    .m7_rty_o(m7s15_rty),
    .m7_sel_i(m7s15_sel),
    .m7_stb_i(m7s15_stb),
    .m7_we_i(m7s15_we),
    .rst_i(_0082_),
    .wb_ack_i(i_s15_ack_i),
    .wb_addr_o(i_s15_addr_o),
    .wb_cyc_o(i_s15_cyc_o),
    .wb_data_i(i_s15_data_i),
    .wb_data_o(i_s15_data_o),
    .wb_err_i(i_s15_err_i),
    .wb_rty_i(i_s15_rty_i),
    .wb_sel_o(i_s15_sel_o),
    .wb_stb_o(i_s15_stb_o),
    .wb_we_o(i_s15_we_o)
  );
\$paramod$babc7f28591f52523637895ab98a5c04b5a93873\wb_conmax_slave_if   s2 (
    .clk_i(_0001_),
    .conf(conf2),
    .m0_ack_o(m0s2_ack),
    .m0_addr_i(m0s2_addr),
    .m0_cyc_i(m0s2_cyc),
    .m0_data_i(m0s2_data_o),
    .m0_data_o(m0s2_data_i),
    .m0_err_o(m0s2_err),
    .m0_rty_o(m0s2_rty),
    .m0_sel_i(m0s2_sel),
    .m0_stb_i(m0s2_stb),
    .m0_we_i(m0s2_we),
    .m1_ack_o(m1s2_ack),
    .m1_addr_i(m1s2_addr),
    .m1_cyc_i(m1s2_cyc),
    .m1_data_i(m1s2_data_o),
    .m1_data_o(m1s2_data_i),
    .m1_err_o(m1s2_err),
    .m1_rty_o(m1s2_rty),
    .m1_sel_i(m1s2_sel),
    .m1_stb_i(m1s2_stb),
    .m1_we_i(m1s2_we),
    .m2_ack_o(m2s2_ack),
    .m2_addr_i(m2s2_addr),
    .m2_cyc_i(m2s2_cyc),
    .m2_data_i(m2s2_data_o),
    .m2_data_o(m2s2_data_i),
    .m2_err_o(m2s2_err),
    .m2_rty_o(m2s2_rty),
    .m2_sel_i(m2s2_sel),
    .m2_stb_i(m2s2_stb),
    .m2_we_i(m2s2_we),
    .m3_ack_o(m3s2_ack),
    .m3_addr_i(m3s2_addr),
    .m3_cyc_i(m3s2_cyc),
    .m3_data_i(m3s2_data_o),
    .m3_data_o(m3s2_data_i),
    .m3_err_o(m3s2_err),
    .m3_rty_o(m3s2_rty),
    .m3_sel_i(m3s2_sel),
    .m3_stb_i(m3s2_stb),
    .m3_we_i(m3s2_we),
    .m4_ack_o(m4s2_ack),
    .m4_addr_i(m4s2_addr),
    .m4_cyc_i(m4s2_cyc),
    .m4_data_i(m4s2_data_o),
    .m4_data_o(m4s2_data_i),
    .m4_err_o(m4s2_err),
    .m4_rty_o(m4s2_rty),
    .m4_sel_i(m4s2_sel),
    .m4_stb_i(m4s2_stb),
    .m4_we_i(m4s2_we),
    .m5_ack_o(m5s2_ack),
    .m5_addr_i(m5s2_addr),
    .m5_cyc_i(m5s2_cyc),
    .m5_data_i(m5s2_data_o),
    .m5_data_o(m5s2_data_i),
    .m5_err_o(m5s2_err),
    .m5_rty_o(m5s2_rty),
    .m5_sel_i(m5s2_sel),
    .m5_stb_i(m5s2_stb),
    .m5_we_i(m5s2_we),
    .m6_ack_o(m6s2_ack),
    .m6_addr_i(m6s2_addr),
    .m6_cyc_i(m6s2_cyc),
    .m6_data_i(m6s2_data_o),
    .m6_data_o(m6s2_data_i),
    .m6_err_o(m6s2_err),
    .m6_rty_o(m6s2_rty),
    .m6_sel_i(m6s2_sel),
    .m6_stb_i(m6s2_stb),
    .m6_we_i(m6s2_we),
    .m7_ack_o(m7s2_ack),
    .m7_addr_i(m7s2_addr),
    .m7_cyc_i(m7s2_cyc),
    .m7_data_i(m7s2_data_o),
    .m7_data_o(m7s2_data_i),
    .m7_err_o(m7s2_err),
    .m7_rty_o(m7s2_rty),
    .m7_sel_i(m7s2_sel),
    .m7_stb_i(m7s2_stb),
    .m7_we_i(m7s2_we),
    .rst_i(_0082_),
    .wb_ack_i(_0163_),
    .wb_addr_o(_0164_),
    .wb_cyc_o(_0165_),
    .wb_data_i(_0166_),
    .wb_data_o(_0167_),
    .wb_err_i(_0168_),
    .wb_rty_i(_0169_),
    .wb_sel_o(_0170_),
    .wb_stb_o(_0171_),
    .wb_we_o(_0172_)
  );
\$paramod$babc7f28591f52523637895ab98a5c04b5a93873\wb_conmax_slave_if   s3 (
    .clk_i(_0001_),
    .conf(conf3),
    .m0_ack_o(m0s3_ack),
    .m0_addr_i(m0s3_addr),
    .m0_cyc_i(m0s3_cyc),
    .m0_data_i(m0s3_data_o),
    .m0_data_o(m0s3_data_i),
    .m0_err_o(m0s3_err),
    .m0_rty_o(m0s3_rty),
    .m0_sel_i(m0s3_sel),
    .m0_stb_i(m0s3_stb),
    .m0_we_i(m0s3_we),
    .m1_ack_o(m1s3_ack),
    .m1_addr_i(m1s3_addr),
    .m1_cyc_i(m1s3_cyc),
    .m1_data_i(m1s3_data_o),
    .m1_data_o(m1s3_data_i),
    .m1_err_o(m1s3_err),
    .m1_rty_o(m1s3_rty),
    .m1_sel_i(m1s3_sel),
    .m1_stb_i(m1s3_stb),
    .m1_we_i(m1s3_we),
    .m2_ack_o(m2s3_ack),
    .m2_addr_i(m2s3_addr),
    .m2_cyc_i(m2s3_cyc),
    .m2_data_i(m2s3_data_o),
    .m2_data_o(m2s3_data_i),
    .m2_err_o(m2s3_err),
    .m2_rty_o(m2s3_rty),
    .m2_sel_i(m2s3_sel),
    .m2_stb_i(m2s3_stb),
    .m2_we_i(m2s3_we),
    .m3_ack_o(m3s3_ack),
    .m3_addr_i(m3s3_addr),
    .m3_cyc_i(m3s3_cyc),
    .m3_data_i(m3s3_data_o),
    .m3_data_o(m3s3_data_i),
    .m3_err_o(m3s3_err),
    .m3_rty_o(m3s3_rty),
    .m3_sel_i(m3s3_sel),
    .m3_stb_i(m3s3_stb),
    .m3_we_i(m3s3_we),
    .m4_ack_o(m4s3_ack),
    .m4_addr_i(m4s3_addr),
    .m4_cyc_i(m4s3_cyc),
    .m4_data_i(m4s3_data_o),
    .m4_data_o(m4s3_data_i),
    .m4_err_o(m4s3_err),
    .m4_rty_o(m4s3_rty),
    .m4_sel_i(m4s3_sel),
    .m4_stb_i(m4s3_stb),
    .m4_we_i(m4s3_we),
    .m5_ack_o(m5s3_ack),
    .m5_addr_i(m5s3_addr),
    .m5_cyc_i(m5s3_cyc),
    .m5_data_i(m5s3_data_o),
    .m5_data_o(m5s3_data_i),
    .m5_err_o(m5s3_err),
    .m5_rty_o(m5s3_rty),
    .m5_sel_i(m5s3_sel),
    .m5_stb_i(m5s3_stb),
    .m5_we_i(m5s3_we),
    .m6_ack_o(m6s3_ack),
    .m6_addr_i(m6s3_addr),
    .m6_cyc_i(m6s3_cyc),
    .m6_data_i(m6s3_data_o),
    .m6_data_o(m6s3_data_i),
    .m6_err_o(m6s3_err),
    .m6_rty_o(m6s3_rty),
    .m6_sel_i(m6s3_sel),
    .m6_stb_i(m6s3_stb),
    .m6_we_i(m6s3_we),
    .m7_ack_o(m7s3_ack),
    .m7_addr_i(m7s3_addr),
    .m7_cyc_i(m7s3_cyc),
    .m7_data_i(m7s3_data_o),
    .m7_data_o(m7s3_data_i),
    .m7_err_o(m7s3_err),
    .m7_rty_o(m7s3_rty),
    .m7_sel_i(m7s3_sel),
    .m7_stb_i(m7s3_stb),
    .m7_we_i(m7s3_we),
    .rst_i(_0082_),
    .wb_ack_i(_0173_),
    .wb_addr_o(_0174_),
    .wb_cyc_o(_0175_),
    .wb_data_i(_0176_),
    .wb_data_o(_0177_),
    .wb_err_i(_0178_),
    .wb_rty_i(_0179_),
    .wb_sel_o(_0180_),
    .wb_stb_o(_0181_),
    .wb_we_o(_0182_)
  );
\$paramod$babc7f28591f52523637895ab98a5c04b5a93873\wb_conmax_slave_if   s4 (
    .clk_i(_0001_),
    .conf(conf4),
    .m0_ack_o(m0s4_ack),
    .m0_addr_i(m0s4_addr),
    .m0_cyc_i(m0s4_cyc),
    .m0_data_i(m0s4_data_o),
    .m0_data_o(m0s4_data_i),
    .m0_err_o(m0s4_err),
    .m0_rty_o(m0s4_rty),
    .m0_sel_i(m0s4_sel),
    .m0_stb_i(m0s4_stb),
    .m0_we_i(m0s4_we),
    .m1_ack_o(m1s4_ack),
    .m1_addr_i(m1s4_addr),
    .m1_cyc_i(m1s4_cyc),
    .m1_data_i(m1s4_data_o),
    .m1_data_o(m1s4_data_i),
    .m1_err_o(m1s4_err),
    .m1_rty_o(m1s4_rty),
    .m1_sel_i(m1s4_sel),
    .m1_stb_i(m1s4_stb),
    .m1_we_i(m1s4_we),
    .m2_ack_o(m2s4_ack),
    .m2_addr_i(m2s4_addr),
    .m2_cyc_i(m2s4_cyc),
    .m2_data_i(m2s4_data_o),
    .m2_data_o(m2s4_data_i),
    .m2_err_o(m2s4_err),
    .m2_rty_o(m2s4_rty),
    .m2_sel_i(m2s4_sel),
    .m2_stb_i(m2s4_stb),
    .m2_we_i(m2s4_we),
    .m3_ack_o(m3s4_ack),
    .m3_addr_i(m3s4_addr),
    .m3_cyc_i(m3s4_cyc),
    .m3_data_i(m3s4_data_o),
    .m3_data_o(m3s4_data_i),
    .m3_err_o(m3s4_err),
    .m3_rty_o(m3s4_rty),
    .m3_sel_i(m3s4_sel),
    .m3_stb_i(m3s4_stb),
    .m3_we_i(m3s4_we),
    .m4_ack_o(m4s4_ack),
    .m4_addr_i(m4s4_addr),
    .m4_cyc_i(m4s4_cyc),
    .m4_data_i(m4s4_data_o),
    .m4_data_o(m4s4_data_i),
    .m4_err_o(m4s4_err),
    .m4_rty_o(m4s4_rty),
    .m4_sel_i(m4s4_sel),
    .m4_stb_i(m4s4_stb),
    .m4_we_i(m4s4_we),
    .m5_ack_o(m5s4_ack),
    .m5_addr_i(m5s4_addr),
    .m5_cyc_i(m5s4_cyc),
    .m5_data_i(m5s4_data_o),
    .m5_data_o(m5s4_data_i),
    .m5_err_o(m5s4_err),
    .m5_rty_o(m5s4_rty),
    .m5_sel_i(m5s4_sel),
    .m5_stb_i(m5s4_stb),
    .m5_we_i(m5s4_we),
    .m6_ack_o(m6s4_ack),
    .m6_addr_i(m6s4_addr),
    .m6_cyc_i(m6s4_cyc),
    .m6_data_i(m6s4_data_o),
    .m6_data_o(m6s4_data_i),
    .m6_err_o(m6s4_err),
    .m6_rty_o(m6s4_rty),
    .m6_sel_i(m6s4_sel),
    .m6_stb_i(m6s4_stb),
    .m6_we_i(m6s4_we),
    .m7_ack_o(m7s4_ack),
    .m7_addr_i(m7s4_addr),
    .m7_cyc_i(m7s4_cyc),
    .m7_data_i(m7s4_data_o),
    .m7_data_o(m7s4_data_i),
    .m7_err_o(m7s4_err),
    .m7_rty_o(m7s4_rty),
    .m7_sel_i(m7s4_sel),
    .m7_stb_i(m7s4_stb),
    .m7_we_i(m7s4_we),
    .rst_i(_0082_),
    .wb_ack_i(_0183_),
    .wb_addr_o(_0184_),
    .wb_cyc_o(_0185_),
    .wb_data_i(_0186_),
    .wb_data_o(_0187_),
    .wb_err_i(_0188_),
    .wb_rty_i(_0189_),
    .wb_sel_o(_0190_),
    .wb_stb_o(_0191_),
    .wb_we_o(_0192_)
  );
\$paramod$babc7f28591f52523637895ab98a5c04b5a93873\wb_conmax_slave_if   s5 (
    .clk_i(_0001_),
    .conf(conf5),
    .m0_ack_o(m0s5_ack),
    .m0_addr_i(m0s5_addr),
    .m0_cyc_i(m0s5_cyc),
    .m0_data_i(m0s5_data_o),
    .m0_data_o(m0s5_data_i),
    .m0_err_o(m0s5_err),
    .m0_rty_o(m0s5_rty),
    .m0_sel_i(m0s5_sel),
    .m0_stb_i(m0s5_stb),
    .m0_we_i(m0s5_we),
    .m1_ack_o(m1s5_ack),
    .m1_addr_i(m1s5_addr),
    .m1_cyc_i(m1s5_cyc),
    .m1_data_i(m1s5_data_o),
    .m1_data_o(m1s5_data_i),
    .m1_err_o(m1s5_err),
    .m1_rty_o(m1s5_rty),
    .m1_sel_i(m1s5_sel),
    .m1_stb_i(m1s5_stb),
    .m1_we_i(m1s5_we),
    .m2_ack_o(m2s5_ack),
    .m2_addr_i(m2s5_addr),
    .m2_cyc_i(m2s5_cyc),
    .m2_data_i(m2s5_data_o),
    .m2_data_o(m2s5_data_i),
    .m2_err_o(m2s5_err),
    .m2_rty_o(m2s5_rty),
    .m2_sel_i(m2s5_sel),
    .m2_stb_i(m2s5_stb),
    .m2_we_i(m2s5_we),
    .m3_ack_o(m3s5_ack),
    .m3_addr_i(m3s5_addr),
    .m3_cyc_i(m3s5_cyc),
    .m3_data_i(m3s5_data_o),
    .m3_data_o(m3s5_data_i),
    .m3_err_o(m3s5_err),
    .m3_rty_o(m3s5_rty),
    .m3_sel_i(m3s5_sel),
    .m3_stb_i(m3s5_stb),
    .m3_we_i(m3s5_we),
    .m4_ack_o(m4s5_ack),
    .m4_addr_i(m4s5_addr),
    .m4_cyc_i(m4s5_cyc),
    .m4_data_i(m4s5_data_o),
    .m4_data_o(m4s5_data_i),
    .m4_err_o(m4s5_err),
    .m4_rty_o(m4s5_rty),
    .m4_sel_i(m4s5_sel),
    .m4_stb_i(m4s5_stb),
    .m4_we_i(m4s5_we),
    .m5_ack_o(m5s5_ack),
    .m5_addr_i(m5s5_addr),
    .m5_cyc_i(m5s5_cyc),
    .m5_data_i(m5s5_data_o),
    .m5_data_o(m5s5_data_i),
    .m5_err_o(m5s5_err),
    .m5_rty_o(m5s5_rty),
    .m5_sel_i(m5s5_sel),
    .m5_stb_i(m5s5_stb),
    .m5_we_i(m5s5_we),
    .m6_ack_o(m6s5_ack),
    .m6_addr_i(m6s5_addr),
    .m6_cyc_i(m6s5_cyc),
    .m6_data_i(m6s5_data_o),
    .m6_data_o(m6s5_data_i),
    .m6_err_o(m6s5_err),
    .m6_rty_o(m6s5_rty),
    .m6_sel_i(m6s5_sel),
    .m6_stb_i(m6s5_stb),
    .m6_we_i(m6s5_we),
    .m7_ack_o(m7s5_ack),
    .m7_addr_i(m7s5_addr),
    .m7_cyc_i(m7s5_cyc),
    .m7_data_i(m7s5_data_o),
    .m7_data_o(m7s5_data_i),
    .m7_err_o(m7s5_err),
    .m7_rty_o(m7s5_rty),
    .m7_sel_i(m7s5_sel),
    .m7_stb_i(m7s5_stb),
    .m7_we_i(m7s5_we),
    .rst_i(_0082_),
    .wb_ack_i(_0193_),
    .wb_addr_o(_0194_),
    .wb_cyc_o(_0195_),
    .wb_data_i(_0196_),
    .wb_data_o(_0197_),
    .wb_err_i(_0198_),
    .wb_rty_i(_0199_),
    .wb_sel_o(_0200_),
    .wb_stb_o(_0201_),
    .wb_we_o(_0202_)
  );
\$paramod$babc7f28591f52523637895ab98a5c04b5a93873\wb_conmax_slave_if   s6 (
    .clk_i(_0001_),
    .conf(conf6),
    .m0_ack_o(m0s6_ack),
    .m0_addr_i(m0s6_addr),
    .m0_cyc_i(m0s6_cyc),
    .m0_data_i(m0s6_data_o),
    .m0_data_o(m0s6_data_i),
    .m0_err_o(m0s6_err),
    .m0_rty_o(m0s6_rty),
    .m0_sel_i(m0s6_sel),
    .m0_stb_i(m0s6_stb),
    .m0_we_i(m0s6_we),
    .m1_ack_o(m1s6_ack),
    .m1_addr_i(m1s6_addr),
    .m1_cyc_i(m1s6_cyc),
    .m1_data_i(m1s6_data_o),
    .m1_data_o(m1s6_data_i),
    .m1_err_o(m1s6_err),
    .m1_rty_o(m1s6_rty),
    .m1_sel_i(m1s6_sel),
    .m1_stb_i(m1s6_stb),
    .m1_we_i(m1s6_we),
    .m2_ack_o(m2s6_ack),
    .m2_addr_i(m2s6_addr),
    .m2_cyc_i(m2s6_cyc),
    .m2_data_i(m2s6_data_o),
    .m2_data_o(m2s6_data_i),
    .m2_err_o(m2s6_err),
    .m2_rty_o(m2s6_rty),
    .m2_sel_i(m2s6_sel),
    .m2_stb_i(m2s6_stb),
    .m2_we_i(m2s6_we),
    .m3_ack_o(m3s6_ack),
    .m3_addr_i(m3s6_addr),
    .m3_cyc_i(m3s6_cyc),
    .m3_data_i(m3s6_data_o),
    .m3_data_o(m3s6_data_i),
    .m3_err_o(m3s6_err),
    .m3_rty_o(m3s6_rty),
    .m3_sel_i(m3s6_sel),
    .m3_stb_i(m3s6_stb),
    .m3_we_i(m3s6_we),
    .m4_ack_o(m4s6_ack),
    .m4_addr_i(m4s6_addr),
    .m4_cyc_i(m4s6_cyc),
    .m4_data_i(m4s6_data_o),
    .m4_data_o(m4s6_data_i),
    .m4_err_o(m4s6_err),
    .m4_rty_o(m4s6_rty),
    .m4_sel_i(m4s6_sel),
    .m4_stb_i(m4s6_stb),
    .m4_we_i(m4s6_we),
    .m5_ack_o(m5s6_ack),
    .m5_addr_i(m5s6_addr),
    .m5_cyc_i(m5s6_cyc),
    .m5_data_i(m5s6_data_o),
    .m5_data_o(m5s6_data_i),
    .m5_err_o(m5s6_err),
    .m5_rty_o(m5s6_rty),
    .m5_sel_i(m5s6_sel),
    .m5_stb_i(m5s6_stb),
    .m5_we_i(m5s6_we),
    .m6_ack_o(m6s6_ack),
    .m6_addr_i(m6s6_addr),
    .m6_cyc_i(m6s6_cyc),
    .m6_data_i(m6s6_data_o),
    .m6_data_o(m6s6_data_i),
    .m6_err_o(m6s6_err),
    .m6_rty_o(m6s6_rty),
    .m6_sel_i(m6s6_sel),
    .m6_stb_i(m6s6_stb),
    .m6_we_i(m6s6_we),
    .m7_ack_o(m7s6_ack),
    .m7_addr_i(m7s6_addr),
    .m7_cyc_i(m7s6_cyc),
    .m7_data_i(m7s6_data_o),
    .m7_data_o(m7s6_data_i),
    .m7_err_o(m7s6_err),
    .m7_rty_o(m7s6_rty),
    .m7_sel_i(m7s6_sel),
    .m7_stb_i(m7s6_stb),
    .m7_we_i(m7s6_we),
    .rst_i(_0082_),
    .wb_ack_i(_0203_),
    .wb_addr_o(_0204_),
    .wb_cyc_o(_0205_),
    .wb_data_i(_0206_),
    .wb_data_o(_0207_),
    .wb_err_i(_0208_),
    .wb_rty_i(_0209_),
    .wb_sel_o(_0210_),
    .wb_stb_o(_0211_),
    .wb_we_o(_0212_)
  );
\$paramod$babc7f28591f52523637895ab98a5c04b5a93873\wb_conmax_slave_if   s7 (
    .clk_i(_0001_),
    .conf(conf7),
    .m0_ack_o(m0s7_ack),
    .m0_addr_i(m0s7_addr),
    .m0_cyc_i(m0s7_cyc),
    .m0_data_i(m0s7_data_o),
    .m0_data_o(m0s7_data_i),
    .m0_err_o(m0s7_err),
    .m0_rty_o(m0s7_rty),
    .m0_sel_i(m0s7_sel),
    .m0_stb_i(m0s7_stb),
    .m0_we_i(m0s7_we),
    .m1_ack_o(m1s7_ack),
    .m1_addr_i(m1s7_addr),
    .m1_cyc_i(m1s7_cyc),
    .m1_data_i(m1s7_data_o),
    .m1_data_o(m1s7_data_i),
    .m1_err_o(m1s7_err),
    .m1_rty_o(m1s7_rty),
    .m1_sel_i(m1s7_sel),
    .m1_stb_i(m1s7_stb),
    .m1_we_i(m1s7_we),
    .m2_ack_o(m2s7_ack),
    .m2_addr_i(m2s7_addr),
    .m2_cyc_i(m2s7_cyc),
    .m2_data_i(m2s7_data_o),
    .m2_data_o(m2s7_data_i),
    .m2_err_o(m2s7_err),
    .m2_rty_o(m2s7_rty),
    .m2_sel_i(m2s7_sel),
    .m2_stb_i(m2s7_stb),
    .m2_we_i(m2s7_we),
    .m3_ack_o(m3s7_ack),
    .m3_addr_i(m3s7_addr),
    .m3_cyc_i(m3s7_cyc),
    .m3_data_i(m3s7_data_o),
    .m3_data_o(m3s7_data_i),
    .m3_err_o(m3s7_err),
    .m3_rty_o(m3s7_rty),
    .m3_sel_i(m3s7_sel),
    .m3_stb_i(m3s7_stb),
    .m3_we_i(m3s7_we),
    .m4_ack_o(m4s7_ack),
    .m4_addr_i(m4s7_addr),
    .m4_cyc_i(m4s7_cyc),
    .m4_data_i(m4s7_data_o),
    .m4_data_o(m4s7_data_i),
    .m4_err_o(m4s7_err),
    .m4_rty_o(m4s7_rty),
    .m4_sel_i(m4s7_sel),
    .m4_stb_i(m4s7_stb),
    .m4_we_i(m4s7_we),
    .m5_ack_o(m5s7_ack),
    .m5_addr_i(m5s7_addr),
    .m5_cyc_i(m5s7_cyc),
    .m5_data_i(m5s7_data_o),
    .m5_data_o(m5s7_data_i),
    .m5_err_o(m5s7_err),
    .m5_rty_o(m5s7_rty),
    .m5_sel_i(m5s7_sel),
    .m5_stb_i(m5s7_stb),
    .m5_we_i(m5s7_we),
    .m6_ack_o(m6s7_ack),
    .m6_addr_i(m6s7_addr),
    .m6_cyc_i(m6s7_cyc),
    .m6_data_i(m6s7_data_o),
    .m6_data_o(m6s7_data_i),
    .m6_err_o(m6s7_err),
    .m6_rty_o(m6s7_rty),
    .m6_sel_i(m6s7_sel),
    .m6_stb_i(m6s7_stb),
    .m6_we_i(m6s7_we),
    .m7_ack_o(m7s7_ack),
    .m7_addr_i(m7s7_addr),
    .m7_cyc_i(m7s7_cyc),
    .m7_data_i(m7s7_data_o),
    .m7_data_o(m7s7_data_i),
    .m7_err_o(m7s7_err),
    .m7_rty_o(m7s7_rty),
    .m7_sel_i(m7s7_sel),
    .m7_stb_i(m7s7_stb),
    .m7_we_i(m7s7_we),
    .rst_i(_0082_),
    .wb_ack_i(_0213_),
    .wb_addr_o(_0214_),
    .wb_cyc_o(_0215_),
    .wb_data_i(_0216_),
    .wb_data_o(_0217_),
    .wb_err_i(_0218_),
    .wb_rty_i(_0219_),
    .wb_sel_o(_0220_),
    .wb_stb_o(_0221_),
    .wb_we_o(_0222_)
  );
\$paramod$babc7f28591f52523637895ab98a5c04b5a93873\wb_conmax_slave_if   s8 (
    .clk_i(_0001_),
    .conf(conf8),
    .m0_ack_o(m0s8_ack),
    .m0_addr_i(m0s8_addr),
    .m0_cyc_i(m0s8_cyc),
    .m0_data_i(m0s8_data_o),
    .m0_data_o(m0s8_data_i),
    .m0_err_o(m0s8_err),
    .m0_rty_o(m0s8_rty),
    .m0_sel_i(m0s8_sel),
    .m0_stb_i(m0s8_stb),
    .m0_we_i(m0s8_we),
    .m1_ack_o(m1s8_ack),
    .m1_addr_i(m1s8_addr),
    .m1_cyc_i(m1s8_cyc),
    .m1_data_i(m1s8_data_o),
    .m1_data_o(m1s8_data_i),
    .m1_err_o(m1s8_err),
    .m1_rty_o(m1s8_rty),
    .m1_sel_i(m1s8_sel),
    .m1_stb_i(m1s8_stb),
    .m1_we_i(m1s8_we),
    .m2_ack_o(m2s8_ack),
    .m2_addr_i(m2s8_addr),
    .m2_cyc_i(m2s8_cyc),
    .m2_data_i(m2s8_data_o),
    .m2_data_o(m2s8_data_i),
    .m2_err_o(m2s8_err),
    .m2_rty_o(m2s8_rty),
    .m2_sel_i(m2s8_sel),
    .m2_stb_i(m2s8_stb),
    .m2_we_i(m2s8_we),
    .m3_ack_o(m3s8_ack),
    .m3_addr_i(m3s8_addr),
    .m3_cyc_i(m3s8_cyc),
    .m3_data_i(m3s8_data_o),
    .m3_data_o(m3s8_data_i),
    .m3_err_o(m3s8_err),
    .m3_rty_o(m3s8_rty),
    .m3_sel_i(m3s8_sel),
    .m3_stb_i(m3s8_stb),
    .m3_we_i(m3s8_we),
    .m4_ack_o(m4s8_ack),
    .m4_addr_i(m4s8_addr),
    .m4_cyc_i(m4s8_cyc),
    .m4_data_i(m4s8_data_o),
    .m4_data_o(m4s8_data_i),
    .m4_err_o(m4s8_err),
    .m4_rty_o(m4s8_rty),
    .m4_sel_i(m4s8_sel),
    .m4_stb_i(m4s8_stb),
    .m4_we_i(m4s8_we),
    .m5_ack_o(m5s8_ack),
    .m5_addr_i(m5s8_addr),
    .m5_cyc_i(m5s8_cyc),
    .m5_data_i(m5s8_data_o),
    .m5_data_o(m5s8_data_i),
    .m5_err_o(m5s8_err),
    .m5_rty_o(m5s8_rty),
    .m5_sel_i(m5s8_sel),
    .m5_stb_i(m5s8_stb),
    .m5_we_i(m5s8_we),
    .m6_ack_o(m6s8_ack),
    .m6_addr_i(m6s8_addr),
    .m6_cyc_i(m6s8_cyc),
    .m6_data_i(m6s8_data_o),
    .m6_data_o(m6s8_data_i),
    .m6_err_o(m6s8_err),
    .m6_rty_o(m6s8_rty),
    .m6_sel_i(m6s8_sel),
    .m6_stb_i(m6s8_stb),
    .m6_we_i(m6s8_we),
    .m7_ack_o(m7s8_ack),
    .m7_addr_i(m7s8_addr),
    .m7_cyc_i(m7s8_cyc),
    .m7_data_i(m7s8_data_o),
    .m7_data_o(m7s8_data_i),
    .m7_err_o(m7s8_err),
    .m7_rty_o(m7s8_rty),
    .m7_sel_i(m7s8_sel),
    .m7_stb_i(m7s8_stb),
    .m7_we_i(m7s8_we),
    .rst_i(_0082_),
    .wb_ack_i(_0223_),
    .wb_addr_o(_0224_),
    .wb_cyc_o(_0225_),
    .wb_data_i(_0226_),
    .wb_data_o(_0227_),
    .wb_err_i(_0228_),
    .wb_rty_i(_0229_),
    .wb_sel_o(_0230_),
    .wb_stb_o(_0231_),
    .wb_we_o(_0232_)
  );
\$paramod$babc7f28591f52523637895ab98a5c04b5a93873\wb_conmax_slave_if   s9 (
    .clk_i(_0001_),
    .conf(conf9),
    .m0_ack_o(m0s9_ack),
    .m0_addr_i(m0s9_addr),
    .m0_cyc_i(m0s9_cyc),
    .m0_data_i(m0s9_data_o),
    .m0_data_o(m0s9_data_i),
    .m0_err_o(m0s9_err),
    .m0_rty_o(m0s9_rty),
    .m0_sel_i(m0s9_sel),
    .m0_stb_i(m0s9_stb),
    .m0_we_i(m0s9_we),
    .m1_ack_o(m1s9_ack),
    .m1_addr_i(m1s9_addr),
    .m1_cyc_i(m1s9_cyc),
    .m1_data_i(m1s9_data_o),
    .m1_data_o(m1s9_data_i),
    .m1_err_o(m1s9_err),
    .m1_rty_o(m1s9_rty),
    .m1_sel_i(m1s9_sel),
    .m1_stb_i(m1s9_stb),
    .m1_we_i(m1s9_we),
    .m2_ack_o(m2s9_ack),
    .m2_addr_i(m2s9_addr),
    .m2_cyc_i(m2s9_cyc),
    .m2_data_i(m2s9_data_o),
    .m2_data_o(m2s9_data_i),
    .m2_err_o(m2s9_err),
    .m2_rty_o(m2s9_rty),
    .m2_sel_i(m2s9_sel),
    .m2_stb_i(m2s9_stb),
    .m2_we_i(m2s9_we),
    .m3_ack_o(m3s9_ack),
    .m3_addr_i(m3s9_addr),
    .m3_cyc_i(m3s9_cyc),
    .m3_data_i(m3s9_data_o),
    .m3_data_o(m3s9_data_i),
    .m3_err_o(m3s9_err),
    .m3_rty_o(m3s9_rty),
    .m3_sel_i(m3s9_sel),
    .m3_stb_i(m3s9_stb),
    .m3_we_i(m3s9_we),
    .m4_ack_o(m4s9_ack),
    .m4_addr_i(m4s9_addr),
    .m4_cyc_i(m4s9_cyc),
    .m4_data_i(m4s9_data_o),
    .m4_data_o(m4s9_data_i),
    .m4_err_o(m4s9_err),
    .m4_rty_o(m4s9_rty),
    .m4_sel_i(m4s9_sel),
    .m4_stb_i(m4s9_stb),
    .m4_we_i(m4s9_we),
    .m5_ack_o(m5s9_ack),
    .m5_addr_i(m5s9_addr),
    .m5_cyc_i(m5s9_cyc),
    .m5_data_i(m5s9_data_o),
    .m5_data_o(m5s9_data_i),
    .m5_err_o(m5s9_err),
    .m5_rty_o(m5s9_rty),
    .m5_sel_i(m5s9_sel),
    .m5_stb_i(m5s9_stb),
    .m5_we_i(m5s9_we),
    .m6_ack_o(m6s9_ack),
    .m6_addr_i(m6s9_addr),
    .m6_cyc_i(m6s9_cyc),
    .m6_data_i(m6s9_data_o),
    .m6_data_o(m6s9_data_i),
    .m6_err_o(m6s9_err),
    .m6_rty_o(m6s9_rty),
    .m6_sel_i(m6s9_sel),
    .m6_stb_i(m6s9_stb),
    .m6_we_i(m6s9_we),
    .m7_ack_o(m7s9_ack),
    .m7_addr_i(m7s9_addr),
    .m7_cyc_i(m7s9_cyc),
    .m7_data_i(m7s9_data_o),
    .m7_data_o(m7s9_data_i),
    .m7_err_o(m7s9_err),
    .m7_rty_o(m7s9_rty),
    .m7_sel_i(m7s9_sel),
    .m7_stb_i(m7s9_stb),
    .m7_we_i(m7s9_we),
    .rst_i(_0082_),
    .wb_ack_i(_0233_),
    .wb_addr_o(_0234_),
    .wb_cyc_o(_0235_),
    .wb_data_i(_0236_),
    .wb_data_o(_0237_),
    .wb_err_i(_0238_),
    .wb_rty_i(_0239_),
    .wb_sel_o(_0240_),
    .wb_stb_o(_0241_),
    .wb_we_o(_0242_)
  );
endmodule
