module u_xmit(sys_clk,  sys_rst_l, uart_xmitH, xmitH, xmit_dataH, xmit_doneH);
wire  [4:0] _000_;
wire  [3:0] _001_;
wire  [7:0] _002_;
wire  _003_;
wire  _004_;
wire  _005_;
wire  _006_;
wire  _007_;
wire  _008_;
wire  _009_;
wire  _010_;
wire  _011_;
wire  _012_;
wire  _013_;
wire  _014_;
wire  _015_;
wire  _016_;
wire  _017_;
wire  _018_;
wire  _019_;
wire  _020_;
wire  _021_;
wire  _022_;
wire  _023_;
wire  _024_;
wire  _025_;
wire  _026_;
wire  _027_;
wire  _028_;
wire  _029_;
wire  _030_;
wire  _031_;
wire  [4:0] _032_;
wire  [4:0] _033_;
wire  [4:0] _034_;
wire  [7:0] _035_;
wire  [7:0] _036_;
wire  [3:0] _037_;
wire  [3:0] _038_;
wire  [3:0] _039_;
wire  _040_;
wire  [1:0] _041_;
wire  [5:0] _042_;
wire  [1:0] _043_;
wire  [4:0] bitCell_cntrH;
wire  [3:0] bitCountH;
wire  [2:0] next_state;
wire  [2:0] state;
input  sys_clk;
wire  sys_clk;
input  sys_rst_l;
wire  sys_rst_l;
output  uart_xmitH;
wire  uart_xmitH;
input  xmitH;
wire  xmitH;
wire  [7:0] xmit_ShiftRegH;
input  [7:0] xmit_dataH;
wire  [7:0] xmit_dataH;
output  xmit_doneH;
wire  xmit_doneH;
wire  xmit_doneInH;
LUT4  #(
    .INIT(16'hcf32)
  ) _044_ (
    .I0(xmitH),
    .I1(state[1]),
    .I2(state[0]),
    .I3(state[2]),
    .O(_009_)
  );
LUT6  #(
    .INIT(64'h3f3300000a003b33)
  ) _045_ (
    .I0(state[0]),
    .I1(xmitH),
    .I2(_042_[0]),
    .I3(_042_[1]),
    .I4(state[1]),
    .I5(state[2]),
    .O(_010_)
  );
LUT5  #(
    .INIT(32'd268435456)
  ) _046_ (
    .I0(bitCell_cntrH[4]),
    .I1(bitCell_cntrH[0]),
    .I2(bitCell_cntrH[1]),
    .I3(bitCell_cntrH[2]),
    .I4(bitCell_cntrH[3]),
    .O(_042_[1])
  );
LUT4  #(
    .INIT(16'h0100)
  ) _047_ (
    .I0(bitCountH[0]),
    .I1(bitCountH[1]),
    .I2(bitCountH[2]),
    .I3(bitCountH[3]),
    .O(_042_[0])
  );
LUT2  #(
    .INIT(4'h4)
  ) _048_ (
    .I0(_043_[0]),
    .I1(_039_[0]),
    .O(_001_[0])
  );
LUT3  #(
    .INIT(8'h41)
  ) _049_ (
    .I0(xmitH),
    .I1(state[2]),
    .I2(state[1]),
    .O(_043_[0])
  );
LUT2  #(
    .INIT(4'h4)
  ) _050_ (
    .I0(_043_[0]),
    .I1(_039_[1]),
    .O(_001_[1])
  );
LUT2  #(
    .INIT(4'h4)
  ) _051_ (
    .I0(_043_[0]),
    .I1(_039_[2]),
    .O(_001_[2])
  );
LUT2  #(
    .INIT(4'h4)
  ) _052_ (
    .I0(_043_[0]),
    .I1(_039_[3]),
    .O(_001_[3])
  );
LUT5  #(
    .INIT(32'd2899102892)
  ) _053_ (
    .I0(xmit_dataH[0]),
    .I1(xmit_ShiftRegH[1]),
    .I2(xmitH),
    .I3(state[1]),
    .I4(state[2]),
    .O(_002_[0])
  );
LUT5  #(
    .INIT(32'd2899102892)
  ) _054_ (
    .I0(xmit_dataH[1]),
    .I1(xmit_ShiftRegH[2]),
    .I2(xmitH),
    .I3(state[1]),
    .I4(state[2]),
    .O(_002_[1])
  );
LUT5  #(
    .INIT(32'd2899102892)
  ) _055_ (
    .I0(xmit_dataH[2]),
    .I1(xmit_ShiftRegH[3]),
    .I2(xmitH),
    .I3(state[1]),
    .I4(state[2]),
    .O(_002_[2])
  );
LUT5  #(
    .INIT(32'd2899102892)
  ) _056_ (
    .I0(xmit_dataH[3]),
    .I1(xmit_ShiftRegH[4]),
    .I2(xmitH),
    .I3(state[1]),
    .I4(state[2]),
    .O(_002_[3])
  );
LUT5  #(
    .INIT(32'd2899102892)
  ) _057_ (
    .I0(xmit_dataH[4]),
    .I1(xmit_ShiftRegH[5]),
    .I2(xmitH),
    .I3(state[1]),
    .I4(state[2]),
    .O(_002_[4])
  );
LUT5  #(
    .INIT(32'd2899102892)
  ) _058_ (
    .I0(xmit_dataH[5]),
    .I1(xmit_ShiftRegH[6]),
    .I2(xmitH),
    .I3(state[1]),
    .I4(state[2]),
    .O(_002_[5])
  );
LUT5  #(
    .INIT(32'd2899102892)
  ) _059_ (
    .I0(xmit_dataH[6]),
    .I1(xmit_ShiftRegH[7]),
    .I2(xmitH),
    .I3(state[1]),
    .I4(state[2]),
    .O(_002_[6])
  );
LUT2  #(
    .INIT(4'h4)
  ) _060_ (
    .I0(_041_[0]),
    .I1(_034_[0]),
    .O(_000_[0])
  );
LUT2  #(
    .INIT(4'h1)
  ) _061_ (
    .I0(state[1]),
    .I1(state[0]),
    .O(_005_)
  );
LUT2  #(
    .INIT(4'h1)
  ) _062_ (
    .I0(state[1]),
    .I1(state[0]),
    .O(_006_)
  );
MUXF7  _063_ (
    .I0(_005_),
    .I1(_006_),
    .O(_003_),
    .S(bitCell_cntrH[2])
  );
LUT2  #(
    .INIT(4'h1)
  ) _064_ (
    .I0(state[1]),
    .I1(state[0]),
    .O(_007_)
  );
LUT6  #(
    .INIT(64'h040b575d00005555)
  ) _065_ (
    .I0(state[1]),
    .I1(state[2]),
    .I2(bitCell_cntrH[4]),
    .I3(bitCell_cntrH[0]),
    .I4(state[0]),
    .I5(bitCell_cntrH[1]),
    .O(_008_)
  );
MUXF7  _066_ (
    .I0(_007_),
    .I1(_008_),
    .O(_004_),
    .S(bitCell_cntrH[2])
  );
MUXF8  _067_ (
    .I0(_003_),
    .I1(_004_),
    .O(_041_[0]),
    .S(bitCell_cntrH[3])
  );
LUT2  #(
    .INIT(4'h4)
  ) _068_ (
    .I0(_041_[0]),
    .I1(_034_[1]),
    .O(_000_[1])
  );
LUT2  #(
    .INIT(4'h4)
  ) _069_ (
    .I0(_041_[0]),
    .I1(_034_[2]),
    .O(_000_[2])
  );
LUT2  #(
    .INIT(4'h4)
  ) _070_ (
    .I0(_041_[0]),
    .I1(_034_[3]),
    .O(_000_[3])
  );
LUT2  #(
    .INIT(4'h4)
  ) _071_ (
    .I0(_041_[0]),
    .I1(_034_[4]),
    .O(_000_[4])
  );
LUT6  #(
    .INIT(64'h00ffffffb0b0f000)
  ) _072_ (
    .I0(_042_[0]),
    .I1(_042_[1]),
    .I2(state[1]),
    .I3(_042_[3]),
    .I4(state[0]),
    .I5(state[2]),
    .O(next_state[0])
  );
LUT5  #(
    .INIT(32'd1073741824)
  ) _073_ (
    .I0(bitCell_cntrH[4]),
    .I1(bitCell_cntrH[0]),
    .I2(bitCell_cntrH[1]),
    .I3(bitCell_cntrH[2]),
    .I4(bitCell_cntrH[3]),
    .O(_042_[3])
  );
LUT5  #(
    .INIT(32'd255791018)
  ) _074_ (
    .I0(xmitH),
    .I1(_042_[1]),
    .I2(state[0]),
    .I3(state[2]),
    .I4(state[1]),
    .O(next_state[1])
  );
LUT5  #(
    .INIT(32'd260571136)
  ) _075_ (
    .I0(_042_[1]),
    .I1(state[1]),
    .I2(_042_[3]),
    .I3(state[2]),
    .I4(state[0]),
    .O(next_state[2])
  );
LUT5  #(
    .INIT(32'd260571151)
  ) _076_ (
    .I0(_042_[3]),
    .I1(state[0]),
    .I2(xmitH),
    .I3(state[1]),
    .I4(state[2]),
    .O(xmit_doneInH)
  );
LUT4  #(
    .INIT(16'h2c0b)
  ) _077_ (
    .I0(xmit_ShiftRegH[0]),
    .I1(state[2]),
    .I2(state[1]),
    .I3(state[0]),
    .O(uart_xmitH)
  );
INV  _078_ (
    .I(sys_rst_l),
    .O(_011_)
  );
INV  _079_ (
    .I(bitCountH[0]),
    .O(_038_[0])
  );
INV  _080_ (
    .I(bitCell_cntrH[0]),
    .O(_033_[0])
  );
INV  _081_ (
    .I(sys_rst_l),
    .O(_012_)
  );
INV  _082_ (
    .I(sys_rst_l),
    .O(_013_)
  );
INV  _083_ (
    .I(sys_rst_l),
    .O(_014_)
  );
INV  _084_ (
    .I(sys_rst_l),
    .O(_015_)
  );
INV  _085_ (
    .I(sys_rst_l),
    .O(_016_)
  );
INV  _086_ (
    .I(sys_rst_l),
    .O(_017_)
  );
INV  _087_ (
    .I(sys_rst_l),
    .O(_018_)
  );
INV  _088_ (
    .I(sys_rst_l),
    .O(_019_)
  );
INV  _089_ (
    .I(sys_rst_l),
    .O(_020_)
  );
INV  _090_ (
    .I(sys_rst_l),
    .O(_021_)
  );
INV  _091_ (
    .I(sys_rst_l),
    .O(_022_)
  );
INV  _092_ (
    .I(sys_rst_l),
    .O(_023_)
  );
INV  _093_ (
    .I(sys_rst_l),
    .O(_024_)
  );
INV  _094_ (
    .I(sys_rst_l),
    .O(_025_)
  );
INV  _095_ (
    .I(sys_rst_l),
    .O(_026_)
  );
INV  _096_ (
    .I(sys_rst_l),
    .O(_027_)
  );
INV  _097_ (
    .I(sys_rst_l),
    .O(_028_)
  );
INV  _098_ (
    .I(sys_rst_l),
    .O(_029_)
  );
INV  _099_ (
    .I(sys_rst_l),
    .O(_030_)
  );
INV  _100_ (
    .I(sys_rst_l),
    .O(_031_)
  );
CARRY4  _101_ (
    .CI(1'h0),
    .CO(_032_[3:0]),
    .CYINIT(1'h0),
    .DI(4'h1),
    .O(_034_[3:0]),
    .S({ bitCell_cntrH[3:1], _033_[0] })
  );
CARRY4  _102_ (
    .CI(_032_[3]),
    .CO({ _035_[7:5], _032_[4] }),
    .CYINIT(1'h0),
    .DI(4'h0),
    .O({ _036_[7:5], _034_[4] }),
    .S({ 3'h0, bitCell_cntrH[4] })
  );
CARRY4  _103_ (
    .CI(1'h0),
    .CO(_037_),
    .CYINIT(1'h0),
    .DI(4'h1),
    .O(_039_),
    .S({ bitCountH[3:1], _038_[0] })
  );
FDCE  #(
    .INIT(1'hx)
  ) _104_ (
    .C(sys_clk),
    .CE(1'h1),
    .CLR(_011_),
    .D(xmit_doneInH),
    .Q(xmit_doneH)
  );
FDCE  #(
    .INIT(1'hx)
  ) _105_ (
    .C(sys_clk),
    .CE(1'h1),
    .CLR(_012_),
    .D(next_state[0]),
    .Q(state[0])
  );
FDCE  #(
    .INIT(1'hx)
  ) _106_ (
    .C(sys_clk),
    .CE(1'h1),
    .CLR(_013_),
    .D(next_state[1]),
    .Q(state[1])
  );
FDCE  #(
    .INIT(1'hx)
  ) _107_ (
    .C(sys_clk),
    .CE(1'h1),
    .CLR(_014_),
    .D(next_state[2]),
    .Q(state[2])
  );
FDCE  #(
    .INIT(1'hx)
  ) _108_ (
    .C(sys_clk),
    .CE(_010_),
    .CLR(_015_),
    .D(_001_[0]),
    .Q(bitCountH[0])
  );
FDCE  #(
    .INIT(1'hx)
  ) _109_ (
    .C(sys_clk),
    .CE(_010_),
    .CLR(_016_),
    .D(_001_[1]),
    .Q(bitCountH[1])
  );
FDCE  #(
    .INIT(1'hx)
  ) _110_ (
    .C(sys_clk),
    .CE(_010_),
    .CLR(_017_),
    .D(_001_[2]),
    .Q(bitCountH[2])
  );
FDCE  #(
    .INIT(1'hx)
  ) _111_ (
    .C(sys_clk),
    .CE(_010_),
    .CLR(_018_),
    .D(_001_[3]),
    .Q(bitCountH[3])
  );
FDCE  #(
    .INIT(1'hx)
  ) _112_ (
    .C(sys_clk),
    .CE(1'h1),
    .CLR(_019_),
    .D(_000_[0]),
    .Q(bitCell_cntrH[0])
  );
FDCE  #(
    .INIT(1'hx)
  ) _113_ (
    .C(sys_clk),
    .CE(1'h1),
    .CLR(_020_),
    .D(_000_[1]),
    .Q(bitCell_cntrH[1])
  );
FDCE  #(
    .INIT(1'hx)
  ) _114_ (
    .C(sys_clk),
    .CE(1'h1),
    .CLR(_021_),
    .D(_000_[2]),
    .Q(bitCell_cntrH[2])
  );
FDCE  #(
    .INIT(1'hx)
  ) _115_ (
    .C(sys_clk),
    .CE(1'h1),
    .CLR(_022_),
    .D(_000_[3]),
    .Q(bitCell_cntrH[3])
  );
FDCE  #(
    .INIT(1'hx)
  ) _116_ (
    .C(sys_clk),
    .CE(1'h1),
    .CLR(_023_),
    .D(_000_[4]),
    .Q(bitCell_cntrH[4])
  );
FDCE  #(
    .INIT(1'hx)
  ) _117_ (
    .C(sys_clk),
    .CE(_009_),
    .CLR(_024_),
    .D(_002_[0]),
    .Q(xmit_ShiftRegH[0])
  );
FDCE  #(
    .INIT(1'hx)
  ) _118_ (
    .C(sys_clk),
    .CE(_009_),
    .CLR(_025_),
    .D(_002_[1]),
    .Q(xmit_ShiftRegH[1])
  );
FDCE  #(
    .INIT(1'hx)
  ) _119_ (
    .C(sys_clk),
    .CE(_009_),
    .CLR(_026_),
    .D(_002_[2]),
    .Q(xmit_ShiftRegH[2])
  );
FDCE  #(
    .INIT(1'hx)
  ) _120_ (
    .C(sys_clk),
    .CE(_009_),
    .CLR(_027_),
    .D(_002_[3]),
    .Q(xmit_ShiftRegH[3])
  );
FDCE  #(
    .INIT(1'hx)
  ) _121_ (
    .C(sys_clk),
    .CE(_009_),
    .CLR(_028_),
    .D(_002_[4]),
    .Q(xmit_ShiftRegH[4])
  );
FDCE  #(
    .INIT(1'hx)
  ) _122_ (
    .C(sys_clk),
    .CE(_009_),
    .CLR(_029_),
    .D(_002_[5]),
    .Q(xmit_ShiftRegH[5])
  );
FDCE  #(
    .INIT(1'hx)
  ) _123_ (
    .C(sys_clk),
    .CE(_009_),
    .CLR(_030_),
    .D(_002_[6]),
    .Q(xmit_ShiftRegH[6])
  );
FDCE  #(
    .INIT(1'hx)
  ) _124_ (
    .C(sys_clk),
    .CE(1'h1),
    .CLR(_031_),
    .D(_040_),
    .Q(xmit_ShiftRegH[7])
  );
LUT6  #(
    .INIT(64'hf0aabbf0ffaabbee)
  ) _125_ (
    .I0(xmit_ShiftRegH[7]),
    .I1(state[0]),
    .I2(xmit_dataH[7]),
    .I3(state[2]),
    .I4(state[1]),
    .I5(xmitH),
    .O(_040_)
  );
assign  { _042_[5:4], _042_[2] } = { state[2], state[0], state[1] };
assign  _043_[1] = _039_[0];
assign  _041_[1] = _034_[1];
assign  _033_[4:1] = bitCell_cntrH[4:1];
assign  _035_[4:0] = _032_;
assign  _036_[4:0] = _034_;
assign  _038_[3:1] = bitCountH[3:1];
endmodule
