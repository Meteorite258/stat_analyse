module AES_Comp_DecCore(di,  ki, Rrg, Kgen, \do , ko);
wire  [7:0] _000_;
wire  _001_;
wire  _002_;
wire  _003_;
wire  _004_;
wire  _005_;
wire  _006_;
wire  _007_;
wire  _008_;
wire  _009_;
wire  _010_;
wire  [6:0] _011_;
wire  _012_;
wire  _013_;
wire  _014_;
wire  [6:0] _015_;
wire  _016_;
wire  _017_;
wire  _018_;
wire  _019_;
wire  _020_;
wire  [6:0] _021_;
wire  _022_;
wire  _023_;
wire  _024_;
wire  [6:0] _025_;
wire  _026_;
wire  _027_;
wire  _028_;
wire  _029_;
wire  _030_;
wire  _031_;
wire  _032_;
wire  _033_;
wire  _034_;
wire  _035_;
wire  _036_;
wire  _037_;
wire  _038_;
wire  _039_;
wire  _040_;
wire  _041_;
wire  _042_;
wire  _043_;
wire  _044_;
wire  _045_;
wire  _046_;
wire  _047_;
wire  _048_;
wire  _049_;
wire  _050_;
wire  _051_;
wire  _052_;
wire  _053_;
wire  _054_;
wire  _055_;
wire  _056_;
wire  _057_;
wire  _058_;
wire  _059_;
wire  _060_;
wire  _061_;
wire  _062_;
wire  _063_;
wire  _064_;
wire  _065_;
wire  _066_;
wire  _067_;
wire  _068_;
wire  _069_;
wire  _070_;
wire  _071_;
wire  _072_;
wire  _073_;
wire  _074_;
wire  _075_;
wire  [5:0] _076_;
wire  [5:0] _077_;
wire  [5:0] _078_;
wire  [5:0] _079_;
wire  [5:0] _080_;
wire  [5:0] _081_;
input  Kgen;
wire  Kgen;
input  [9:0] Rrg;
wire  [9:0] Rrg;
input  [127:0] di;
wire  [127:0] di;
output  [127:0] \do ;
wire  [127:0] \do ;
wire  [127:0] dx;
input  [127:0] ki;
wire  [127:0] ki;
output  [127:0] ko;
wire  [127:0] ko;
wire  [127:0] mx;
wire  [9:0] \rcon$func$AES_Comp.v:408$441.x ;
wire  [9:0] \rcon$func$AES_Comp.v:412$442.x ;
wire  [127:0] sb;
wire  [31:0] so;
wire  [127:0] sr;
LUT3  #(
    .INIT(8'hac)
  ) _082_ (
    .I0(di[0]),
    .I1(mx[0]),
    .I2(Rrg[8]),
    .O(dx[0])
  );
LUT3  #(
    .INIT(8'hca)
  ) _083_ (
    .I0(mx[1]),
    .I1(di[1]),
    .I2(Rrg[8]),
    .O(dx[1])
  );
LUT3  #(
    .INIT(8'hca)
  ) _084_ (
    .I0(mx[2]),
    .I1(di[2]),
    .I2(Rrg[8]),
    .O(dx[2])
  );
LUT3  #(
    .INIT(8'hca)
  ) _085_ (
    .I0(mx[3]),
    .I1(di[3]),
    .I2(Rrg[8]),
    .O(dx[3])
  );
LUT3  #(
    .INIT(8'hca)
  ) _086_ (
    .I0(mx[4]),
    .I1(di[4]),
    .I2(Rrg[8]),
    .O(dx[4])
  );
LUT3  #(
    .INIT(8'hca)
  ) _087_ (
    .I0(mx[5]),
    .I1(di[5]),
    .I2(Rrg[8]),
    .O(dx[5])
  );
LUT3  #(
    .INIT(8'hca)
  ) _088_ (
    .I0(mx[6]),
    .I1(di[6]),
    .I2(Rrg[8]),
    .O(dx[6])
  );
LUT3  #(
    .INIT(8'hca)
  ) _089_ (
    .I0(mx[7]),
    .I1(di[7]),
    .I2(Rrg[8]),
    .O(dx[7])
  );
LUT3  #(
    .INIT(8'hca)
  ) _090_ (
    .I0(mx[8]),
    .I1(di[8]),
    .I2(Rrg[8]),
    .O(dx[8])
  );
LUT3  #(
    .INIT(8'hca)
  ) _091_ (
    .I0(mx[9]),
    .I1(di[9]),
    .I2(Rrg[8]),
    .O(dx[9])
  );
LUT3  #(
    .INIT(8'hca)
  ) _092_ (
    .I0(mx[10]),
    .I1(di[10]),
    .I2(Rrg[8]),
    .O(dx[10])
  );
LUT3  #(
    .INIT(8'hca)
  ) _093_ (
    .I0(mx[11]),
    .I1(di[11]),
    .I2(Rrg[8]),
    .O(dx[11])
  );
LUT3  #(
    .INIT(8'hca)
  ) _094_ (
    .I0(mx[12]),
    .I1(di[12]),
    .I2(Rrg[8]),
    .O(dx[12])
  );
LUT3  #(
    .INIT(8'hca)
  ) _095_ (
    .I0(mx[13]),
    .I1(di[13]),
    .I2(Rrg[8]),
    .O(dx[13])
  );
LUT3  #(
    .INIT(8'hca)
  ) _096_ (
    .I0(mx[14]),
    .I1(di[14]),
    .I2(Rrg[8]),
    .O(dx[14])
  );
LUT3  #(
    .INIT(8'hca)
  ) _097_ (
    .I0(mx[15]),
    .I1(di[15]),
    .I2(Rrg[8]),
    .O(dx[15])
  );
LUT3  #(
    .INIT(8'hca)
  ) _098_ (
    .I0(mx[16]),
    .I1(di[16]),
    .I2(Rrg[8]),
    .O(dx[16])
  );
LUT3  #(
    .INIT(8'hca)
  ) _099_ (
    .I0(mx[17]),
    .I1(di[17]),
    .I2(Rrg[8]),
    .O(dx[17])
  );
LUT3  #(
    .INIT(8'hca)
  ) _100_ (
    .I0(mx[18]),
    .I1(di[18]),
    .I2(Rrg[8]),
    .O(dx[18])
  );
LUT3  #(
    .INIT(8'hca)
  ) _101_ (
    .I0(mx[19]),
    .I1(di[19]),
    .I2(Rrg[8]),
    .O(dx[19])
  );
LUT3  #(
    .INIT(8'hca)
  ) _102_ (
    .I0(mx[20]),
    .I1(di[20]),
    .I2(Rrg[8]),
    .O(dx[20])
  );
LUT3  #(
    .INIT(8'hca)
  ) _103_ (
    .I0(mx[21]),
    .I1(di[21]),
    .I2(Rrg[8]),
    .O(dx[21])
  );
LUT3  #(
    .INIT(8'hca)
  ) _104_ (
    .I0(mx[22]),
    .I1(di[22]),
    .I2(Rrg[8]),
    .O(dx[22])
  );
LUT3  #(
    .INIT(8'hca)
  ) _105_ (
    .I0(mx[23]),
    .I1(di[23]),
    .I2(Rrg[8]),
    .O(dx[23])
  );
LUT3  #(
    .INIT(8'hca)
  ) _106_ (
    .I0(mx[24]),
    .I1(di[24]),
    .I2(Rrg[8]),
    .O(dx[24])
  );
LUT3  #(
    .INIT(8'hca)
  ) _107_ (
    .I0(mx[25]),
    .I1(di[25]),
    .I2(Rrg[8]),
    .O(dx[25])
  );
LUT3  #(
    .INIT(8'hca)
  ) _108_ (
    .I0(mx[26]),
    .I1(di[26]),
    .I2(Rrg[8]),
    .O(dx[26])
  );
LUT3  #(
    .INIT(8'hca)
  ) _109_ (
    .I0(mx[27]),
    .I1(di[27]),
    .I2(Rrg[8]),
    .O(dx[27])
  );
LUT3  #(
    .INIT(8'hca)
  ) _110_ (
    .I0(mx[28]),
    .I1(di[28]),
    .I2(Rrg[8]),
    .O(dx[28])
  );
LUT3  #(
    .INIT(8'hca)
  ) _111_ (
    .I0(mx[29]),
    .I1(di[29]),
    .I2(Rrg[8]),
    .O(dx[29])
  );
LUT3  #(
    .INIT(8'hca)
  ) _112_ (
    .I0(mx[30]),
    .I1(di[30]),
    .I2(Rrg[8]),
    .O(dx[30])
  );
LUT3  #(
    .INIT(8'hca)
  ) _113_ (
    .I0(mx[31]),
    .I1(di[31]),
    .I2(Rrg[8]),
    .O(dx[31])
  );
LUT3  #(
    .INIT(8'hca)
  ) _114_ (
    .I0(mx[32]),
    .I1(di[32]),
    .I2(Rrg[8]),
    .O(dx[32])
  );
LUT3  #(
    .INIT(8'hca)
  ) _115_ (
    .I0(mx[33]),
    .I1(di[33]),
    .I2(Rrg[8]),
    .O(dx[33])
  );
LUT3  #(
    .INIT(8'hca)
  ) _116_ (
    .I0(mx[34]),
    .I1(di[34]),
    .I2(Rrg[8]),
    .O(dx[34])
  );
LUT3  #(
    .INIT(8'hca)
  ) _117_ (
    .I0(mx[35]),
    .I1(di[35]),
    .I2(Rrg[8]),
    .O(dx[35])
  );
LUT3  #(
    .INIT(8'hca)
  ) _118_ (
    .I0(mx[36]),
    .I1(di[36]),
    .I2(Rrg[8]),
    .O(dx[36])
  );
LUT3  #(
    .INIT(8'hca)
  ) _119_ (
    .I0(mx[37]),
    .I1(di[37]),
    .I2(Rrg[8]),
    .O(dx[37])
  );
LUT3  #(
    .INIT(8'hca)
  ) _120_ (
    .I0(mx[38]),
    .I1(di[38]),
    .I2(Rrg[8]),
    .O(dx[38])
  );
LUT3  #(
    .INIT(8'hca)
  ) _121_ (
    .I0(mx[39]),
    .I1(di[39]),
    .I2(Rrg[8]),
    .O(dx[39])
  );
LUT3  #(
    .INIT(8'hca)
  ) _122_ (
    .I0(mx[40]),
    .I1(di[40]),
    .I2(Rrg[8]),
    .O(dx[40])
  );
LUT3  #(
    .INIT(8'hca)
  ) _123_ (
    .I0(mx[41]),
    .I1(di[41]),
    .I2(Rrg[8]),
    .O(dx[41])
  );
LUT3  #(
    .INIT(8'hca)
  ) _124_ (
    .I0(mx[42]),
    .I1(di[42]),
    .I2(Rrg[8]),
    .O(dx[42])
  );
LUT3  #(
    .INIT(8'hca)
  ) _125_ (
    .I0(mx[43]),
    .I1(di[43]),
    .I2(Rrg[8]),
    .O(dx[43])
  );
LUT3  #(
    .INIT(8'hca)
  ) _126_ (
    .I0(mx[44]),
    .I1(di[44]),
    .I2(Rrg[8]),
    .O(dx[44])
  );
LUT3  #(
    .INIT(8'hca)
  ) _127_ (
    .I0(mx[45]),
    .I1(di[45]),
    .I2(Rrg[8]),
    .O(dx[45])
  );
LUT3  #(
    .INIT(8'hca)
  ) _128_ (
    .I0(mx[46]),
    .I1(di[46]),
    .I2(Rrg[8]),
    .O(dx[46])
  );
LUT3  #(
    .INIT(8'hca)
  ) _129_ (
    .I0(mx[47]),
    .I1(di[47]),
    .I2(Rrg[8]),
    .O(dx[47])
  );
LUT3  #(
    .INIT(8'hca)
  ) _130_ (
    .I0(mx[48]),
    .I1(di[48]),
    .I2(Rrg[8]),
    .O(dx[48])
  );
LUT3  #(
    .INIT(8'hca)
  ) _131_ (
    .I0(mx[49]),
    .I1(di[49]),
    .I2(Rrg[8]),
    .O(dx[49])
  );
LUT3  #(
    .INIT(8'hca)
  ) _132_ (
    .I0(mx[50]),
    .I1(di[50]),
    .I2(Rrg[8]),
    .O(dx[50])
  );
LUT3  #(
    .INIT(8'hca)
  ) _133_ (
    .I0(mx[51]),
    .I1(di[51]),
    .I2(Rrg[8]),
    .O(dx[51])
  );
LUT3  #(
    .INIT(8'hca)
  ) _134_ (
    .I0(mx[52]),
    .I1(di[52]),
    .I2(Rrg[8]),
    .O(dx[52])
  );
LUT3  #(
    .INIT(8'hca)
  ) _135_ (
    .I0(mx[53]),
    .I1(di[53]),
    .I2(Rrg[8]),
    .O(dx[53])
  );
LUT3  #(
    .INIT(8'hca)
  ) _136_ (
    .I0(mx[54]),
    .I1(di[54]),
    .I2(Rrg[8]),
    .O(dx[54])
  );
LUT3  #(
    .INIT(8'hca)
  ) _137_ (
    .I0(mx[55]),
    .I1(di[55]),
    .I2(Rrg[8]),
    .O(dx[55])
  );
LUT3  #(
    .INIT(8'hca)
  ) _138_ (
    .I0(mx[56]),
    .I1(di[56]),
    .I2(Rrg[8]),
    .O(dx[56])
  );
LUT3  #(
    .INIT(8'hca)
  ) _139_ (
    .I0(mx[57]),
    .I1(di[57]),
    .I2(Rrg[8]),
    .O(dx[57])
  );
LUT3  #(
    .INIT(8'hca)
  ) _140_ (
    .I0(mx[58]),
    .I1(di[58]),
    .I2(Rrg[8]),
    .O(dx[58])
  );
LUT3  #(
    .INIT(8'hca)
  ) _141_ (
    .I0(mx[59]),
    .I1(di[59]),
    .I2(Rrg[8]),
    .O(dx[59])
  );
LUT3  #(
    .INIT(8'hca)
  ) _142_ (
    .I0(mx[60]),
    .I1(di[60]),
    .I2(Rrg[8]),
    .O(dx[60])
  );
LUT3  #(
    .INIT(8'hca)
  ) _143_ (
    .I0(mx[61]),
    .I1(di[61]),
    .I2(Rrg[8]),
    .O(dx[61])
  );
LUT3  #(
    .INIT(8'hca)
  ) _144_ (
    .I0(mx[62]),
    .I1(di[62]),
    .I2(Rrg[8]),
    .O(dx[62])
  );
LUT3  #(
    .INIT(8'hca)
  ) _145_ (
    .I0(mx[63]),
    .I1(di[63]),
    .I2(Rrg[8]),
    .O(dx[63])
  );
LUT3  #(
    .INIT(8'hca)
  ) _146_ (
    .I0(mx[64]),
    .I1(di[64]),
    .I2(Rrg[8]),
    .O(dx[64])
  );
LUT3  #(
    .INIT(8'hca)
  ) _147_ (
    .I0(mx[65]),
    .I1(di[65]),
    .I2(Rrg[8]),
    .O(dx[65])
  );
LUT3  #(
    .INIT(8'hca)
  ) _148_ (
    .I0(mx[66]),
    .I1(di[66]),
    .I2(Rrg[8]),
    .O(dx[66])
  );
LUT3  #(
    .INIT(8'hca)
  ) _149_ (
    .I0(mx[67]),
    .I1(di[67]),
    .I2(Rrg[8]),
    .O(dx[67])
  );
LUT3  #(
    .INIT(8'hca)
  ) _150_ (
    .I0(mx[68]),
    .I1(di[68]),
    .I2(Rrg[8]),
    .O(dx[68])
  );
LUT3  #(
    .INIT(8'hca)
  ) _151_ (
    .I0(mx[69]),
    .I1(di[69]),
    .I2(Rrg[8]),
    .O(dx[69])
  );
LUT3  #(
    .INIT(8'hca)
  ) _152_ (
    .I0(mx[70]),
    .I1(di[70]),
    .I2(Rrg[8]),
    .O(dx[70])
  );
LUT3  #(
    .INIT(8'hca)
  ) _153_ (
    .I0(mx[71]),
    .I1(di[71]),
    .I2(Rrg[8]),
    .O(dx[71])
  );
LUT3  #(
    .INIT(8'hca)
  ) _154_ (
    .I0(mx[72]),
    .I1(di[72]),
    .I2(Rrg[8]),
    .O(dx[72])
  );
LUT3  #(
    .INIT(8'hca)
  ) _155_ (
    .I0(mx[73]),
    .I1(di[73]),
    .I2(Rrg[8]),
    .O(dx[73])
  );
LUT3  #(
    .INIT(8'hca)
  ) _156_ (
    .I0(mx[74]),
    .I1(di[74]),
    .I2(Rrg[8]),
    .O(dx[74])
  );
LUT3  #(
    .INIT(8'hca)
  ) _157_ (
    .I0(mx[75]),
    .I1(di[75]),
    .I2(Rrg[8]),
    .O(dx[75])
  );
LUT3  #(
    .INIT(8'hca)
  ) _158_ (
    .I0(mx[76]),
    .I1(di[76]),
    .I2(Rrg[8]),
    .O(dx[76])
  );
LUT3  #(
    .INIT(8'hca)
  ) _159_ (
    .I0(mx[77]),
    .I1(di[77]),
    .I2(Rrg[8]),
    .O(dx[77])
  );
LUT3  #(
    .INIT(8'hca)
  ) _160_ (
    .I0(mx[78]),
    .I1(di[78]),
    .I2(Rrg[8]),
    .O(dx[78])
  );
LUT3  #(
    .INIT(8'hca)
  ) _161_ (
    .I0(mx[79]),
    .I1(di[79]),
    .I2(Rrg[8]),
    .O(dx[79])
  );
LUT3  #(
    .INIT(8'hca)
  ) _162_ (
    .I0(mx[80]),
    .I1(di[80]),
    .I2(Rrg[8]),
    .O(dx[80])
  );
LUT3  #(
    .INIT(8'hca)
  ) _163_ (
    .I0(mx[81]),
    .I1(di[81]),
    .I2(Rrg[8]),
    .O(dx[81])
  );
LUT3  #(
    .INIT(8'hca)
  ) _164_ (
    .I0(mx[82]),
    .I1(di[82]),
    .I2(Rrg[8]),
    .O(dx[82])
  );
LUT3  #(
    .INIT(8'hca)
  ) _165_ (
    .I0(mx[83]),
    .I1(di[83]),
    .I2(Rrg[8]),
    .O(dx[83])
  );
LUT3  #(
    .INIT(8'hca)
  ) _166_ (
    .I0(mx[84]),
    .I1(di[84]),
    .I2(Rrg[8]),
    .O(dx[84])
  );
LUT3  #(
    .INIT(8'hca)
  ) _167_ (
    .I0(mx[85]),
    .I1(di[85]),
    .I2(Rrg[8]),
    .O(dx[85])
  );
LUT3  #(
    .INIT(8'hca)
  ) _168_ (
    .I0(mx[86]),
    .I1(di[86]),
    .I2(Rrg[8]),
    .O(dx[86])
  );
LUT3  #(
    .INIT(8'hca)
  ) _169_ (
    .I0(mx[87]),
    .I1(di[87]),
    .I2(Rrg[8]),
    .O(dx[87])
  );
LUT3  #(
    .INIT(8'hca)
  ) _170_ (
    .I0(mx[88]),
    .I1(di[88]),
    .I2(Rrg[8]),
    .O(dx[88])
  );
LUT3  #(
    .INIT(8'hca)
  ) _171_ (
    .I0(mx[89]),
    .I1(di[89]),
    .I2(Rrg[8]),
    .O(dx[89])
  );
LUT3  #(
    .INIT(8'hca)
  ) _172_ (
    .I0(mx[90]),
    .I1(di[90]),
    .I2(Rrg[8]),
    .O(dx[90])
  );
LUT3  #(
    .INIT(8'hca)
  ) _173_ (
    .I0(mx[91]),
    .I1(di[91]),
    .I2(Rrg[8]),
    .O(dx[91])
  );
LUT3  #(
    .INIT(8'hca)
  ) _174_ (
    .I0(mx[92]),
    .I1(di[92]),
    .I2(Rrg[8]),
    .O(dx[92])
  );
LUT3  #(
    .INIT(8'hca)
  ) _175_ (
    .I0(mx[93]),
    .I1(di[93]),
    .I2(Rrg[8]),
    .O(dx[93])
  );
LUT3  #(
    .INIT(8'hca)
  ) _176_ (
    .I0(mx[94]),
    .I1(di[94]),
    .I2(Rrg[8]),
    .O(dx[94])
  );
LUT3  #(
    .INIT(8'hca)
  ) _177_ (
    .I0(mx[95]),
    .I1(di[95]),
    .I2(Rrg[8]),
    .O(dx[95])
  );
LUT3  #(
    .INIT(8'hca)
  ) _178_ (
    .I0(mx[96]),
    .I1(di[96]),
    .I2(Rrg[8]),
    .O(dx[96])
  );
LUT3  #(
    .INIT(8'hca)
  ) _179_ (
    .I0(mx[97]),
    .I1(di[97]),
    .I2(Rrg[8]),
    .O(dx[97])
  );
LUT3  #(
    .INIT(8'hca)
  ) _180_ (
    .I0(mx[98]),
    .I1(di[98]),
    .I2(Rrg[8]),
    .O(dx[98])
  );
LUT3  #(
    .INIT(8'hca)
  ) _181_ (
    .I0(mx[99]),
    .I1(di[99]),
    .I2(Rrg[8]),
    .O(dx[99])
  );
LUT3  #(
    .INIT(8'hca)
  ) _182_ (
    .I0(mx[100]),
    .I1(di[100]),
    .I2(Rrg[8]),
    .O(dx[100])
  );
LUT3  #(
    .INIT(8'hca)
  ) _183_ (
    .I0(mx[101]),
    .I1(di[101]),
    .I2(Rrg[8]),
    .O(dx[101])
  );
LUT3  #(
    .INIT(8'hca)
  ) _184_ (
    .I0(mx[102]),
    .I1(di[102]),
    .I2(Rrg[8]),
    .O(dx[102])
  );
LUT3  #(
    .INIT(8'hca)
  ) _185_ (
    .I0(mx[103]),
    .I1(di[103]),
    .I2(Rrg[8]),
    .O(dx[103])
  );
LUT3  #(
    .INIT(8'hca)
  ) _186_ (
    .I0(mx[104]),
    .I1(di[104]),
    .I2(Rrg[8]),
    .O(dx[104])
  );
LUT3  #(
    .INIT(8'hca)
  ) _187_ (
    .I0(mx[105]),
    .I1(di[105]),
    .I2(Rrg[8]),
    .O(dx[105])
  );
LUT3  #(
    .INIT(8'hca)
  ) _188_ (
    .I0(mx[106]),
    .I1(di[106]),
    .I2(Rrg[8]),
    .O(dx[106])
  );
LUT3  #(
    .INIT(8'hca)
  ) _189_ (
    .I0(mx[107]),
    .I1(di[107]),
    .I2(Rrg[8]),
    .O(dx[107])
  );
LUT3  #(
    .INIT(8'hca)
  ) _190_ (
    .I0(mx[108]),
    .I1(di[108]),
    .I2(Rrg[8]),
    .O(dx[108])
  );
LUT3  #(
    .INIT(8'hca)
  ) _191_ (
    .I0(mx[109]),
    .I1(di[109]),
    .I2(Rrg[8]),
    .O(dx[109])
  );
LUT3  #(
    .INIT(8'hca)
  ) _192_ (
    .I0(mx[110]),
    .I1(di[110]),
    .I2(Rrg[8]),
    .O(dx[110])
  );
LUT3  #(
    .INIT(8'hca)
  ) _193_ (
    .I0(mx[111]),
    .I1(di[111]),
    .I2(Rrg[8]),
    .O(dx[111])
  );
LUT3  #(
    .INIT(8'hca)
  ) _194_ (
    .I0(mx[112]),
    .I1(di[112]),
    .I2(Rrg[8]),
    .O(dx[112])
  );
LUT3  #(
    .INIT(8'hca)
  ) _195_ (
    .I0(mx[113]),
    .I1(di[113]),
    .I2(Rrg[8]),
    .O(dx[113])
  );
LUT3  #(
    .INIT(8'hca)
  ) _196_ (
    .I0(mx[114]),
    .I1(di[114]),
    .I2(Rrg[8]),
    .O(dx[114])
  );
LUT3  #(
    .INIT(8'hca)
  ) _197_ (
    .I0(mx[115]),
    .I1(di[115]),
    .I2(Rrg[8]),
    .O(dx[115])
  );
LUT3  #(
    .INIT(8'hca)
  ) _198_ (
    .I0(mx[116]),
    .I1(di[116]),
    .I2(Rrg[8]),
    .O(dx[116])
  );
LUT3  #(
    .INIT(8'hca)
  ) _199_ (
    .I0(mx[117]),
    .I1(di[117]),
    .I2(Rrg[8]),
    .O(dx[117])
  );
LUT3  #(
    .INIT(8'hca)
  ) _200_ (
    .I0(mx[118]),
    .I1(di[118]),
    .I2(Rrg[8]),
    .O(dx[118])
  );
LUT3  #(
    .INIT(8'hca)
  ) _201_ (
    .I0(mx[119]),
    .I1(di[119]),
    .I2(Rrg[8]),
    .O(dx[119])
  );
LUT3  #(
    .INIT(8'hca)
  ) _202_ (
    .I0(mx[120]),
    .I1(di[120]),
    .I2(Rrg[8]),
    .O(dx[120])
  );
LUT3  #(
    .INIT(8'hca)
  ) _203_ (
    .I0(mx[121]),
    .I1(di[121]),
    .I2(Rrg[8]),
    .O(dx[121])
  );
LUT3  #(
    .INIT(8'hca)
  ) _204_ (
    .I0(mx[122]),
    .I1(di[122]),
    .I2(Rrg[8]),
    .O(dx[122])
  );
LUT3  #(
    .INIT(8'hca)
  ) _205_ (
    .I0(mx[123]),
    .I1(di[123]),
    .I2(Rrg[8]),
    .O(dx[123])
  );
LUT3  #(
    .INIT(8'hca)
  ) _206_ (
    .I0(mx[124]),
    .I1(di[124]),
    .I2(Rrg[8]),
    .O(dx[124])
  );
LUT3  #(
    .INIT(8'hca)
  ) _207_ (
    .I0(mx[125]),
    .I1(di[125]),
    .I2(Rrg[8]),
    .O(dx[125])
  );
LUT3  #(
    .INIT(8'hca)
  ) _208_ (
    .I0(mx[126]),
    .I1(di[126]),
    .I2(Rrg[8]),
    .O(dx[126])
  );
LUT3  #(
    .INIT(8'hca)
  ) _209_ (
    .I0(mx[127]),
    .I1(di[127]),
    .I2(Rrg[8]),
    .O(dx[127])
  );
LUT3  #(
    .INIT(8'hb4)
  ) _210_ (
    .I0(Kgen),
    .I1(ki[56]),
    .I2(ki[24]),
    .O(_044_)
  );
LUT3  #(
    .INIT(8'hb4)
  ) _211_ (
    .I0(Kgen),
    .I1(ki[57]),
    .I2(ki[25]),
    .O(_055_)
  );
LUT3  #(
    .INIT(8'hb4)
  ) _212_ (
    .I0(Kgen),
    .I1(ki[58]),
    .I2(ki[26]),
    .O(_066_)
  );
LUT3  #(
    .INIT(8'hb4)
  ) _213_ (
    .I0(Kgen),
    .I1(ki[59]),
    .I2(ki[27]),
    .O(_069_)
  );
LUT3  #(
    .INIT(8'hb4)
  ) _214_ (
    .I0(Kgen),
    .I1(ki[60]),
    .I2(ki[28]),
    .O(_070_)
  );
LUT3  #(
    .INIT(8'hb4)
  ) _215_ (
    .I0(Kgen),
    .I1(ki[61]),
    .I2(ki[29]),
    .O(_071_)
  );
LUT3  #(
    .INIT(8'hb4)
  ) _216_ (
    .I0(Kgen),
    .I1(ki[62]),
    .I2(ki[30]),
    .O(_072_)
  );
LUT3  #(
    .INIT(8'hb4)
  ) _217_ (
    .I0(Kgen),
    .I1(ki[63]),
    .I2(ki[31]),
    .O(_073_)
  );
LUT3  #(
    .INIT(8'hb4)
  ) _218_ (
    .I0(Kgen),
    .I1(ki[32]),
    .I2(ki[0]),
    .O(_074_)
  );
LUT3  #(
    .INIT(8'hb4)
  ) _219_ (
    .I0(Kgen),
    .I1(ki[33]),
    .I2(ki[1]),
    .O(_075_)
  );
LUT3  #(
    .INIT(8'hb4)
  ) _220_ (
    .I0(Kgen),
    .I1(ki[34]),
    .I2(ki[2]),
    .O(_045_)
  );
LUT3  #(
    .INIT(8'hb4)
  ) _221_ (
    .I0(Kgen),
    .I1(ki[35]),
    .I2(ki[3]),
    .O(_046_)
  );
LUT3  #(
    .INIT(8'hb4)
  ) _222_ (
    .I0(Kgen),
    .I1(ki[36]),
    .I2(ki[4]),
    .O(_047_)
  );
LUT3  #(
    .INIT(8'hb4)
  ) _223_ (
    .I0(Kgen),
    .I1(ki[37]),
    .I2(ki[5]),
    .O(_048_)
  );
LUT3  #(
    .INIT(8'hb4)
  ) _224_ (
    .I0(Kgen),
    .I1(ki[38]),
    .I2(ki[6]),
    .O(_049_)
  );
LUT3  #(
    .INIT(8'hb4)
  ) _225_ (
    .I0(Kgen),
    .I1(ki[39]),
    .I2(ki[7]),
    .O(_050_)
  );
LUT3  #(
    .INIT(8'hb4)
  ) _226_ (
    .I0(Kgen),
    .I1(ki[40]),
    .I2(ki[8]),
    .O(_051_)
  );
LUT3  #(
    .INIT(8'hb4)
  ) _227_ (
    .I0(Kgen),
    .I1(ki[41]),
    .I2(ki[9]),
    .O(_052_)
  );
LUT3  #(
    .INIT(8'hb4)
  ) _228_ (
    .I0(Kgen),
    .I1(ki[42]),
    .I2(ki[10]),
    .O(_053_)
  );
LUT3  #(
    .INIT(8'hb4)
  ) _229_ (
    .I0(Kgen),
    .I1(ki[43]),
    .I2(ki[11]),
    .O(_054_)
  );
LUT3  #(
    .INIT(8'hb4)
  ) _230_ (
    .I0(Kgen),
    .I1(ki[44]),
    .I2(ki[12]),
    .O(_056_)
  );
LUT3  #(
    .INIT(8'hb4)
  ) _231_ (
    .I0(Kgen),
    .I1(ki[45]),
    .I2(ki[13]),
    .O(_057_)
  );
LUT3  #(
    .INIT(8'hb4)
  ) _232_ (
    .I0(Kgen),
    .I1(ki[46]),
    .I2(ki[14]),
    .O(_058_)
  );
LUT3  #(
    .INIT(8'hb4)
  ) _233_ (
    .I0(Kgen),
    .I1(ki[47]),
    .I2(ki[15]),
    .O(_059_)
  );
LUT3  #(
    .INIT(8'hb4)
  ) _234_ (
    .I0(Kgen),
    .I1(ki[48]),
    .I2(ki[16]),
    .O(_060_)
  );
LUT3  #(
    .INIT(8'hb4)
  ) _235_ (
    .I0(Kgen),
    .I1(ki[49]),
    .I2(ki[17]),
    .O(_061_)
  );
LUT3  #(
    .INIT(8'hb4)
  ) _236_ (
    .I0(Kgen),
    .I1(ki[50]),
    .I2(ki[18]),
    .O(_062_)
  );
LUT3  #(
    .INIT(8'hb4)
  ) _237_ (
    .I0(Kgen),
    .I1(ki[51]),
    .I2(ki[19]),
    .O(_063_)
  );
LUT3  #(
    .INIT(8'hb4)
  ) _238_ (
    .I0(Kgen),
    .I1(ki[52]),
    .I2(ki[20]),
    .O(_064_)
  );
LUT3  #(
    .INIT(8'hb4)
  ) _239_ (
    .I0(Kgen),
    .I1(ki[53]),
    .I2(ki[21]),
    .O(_065_)
  );
LUT3  #(
    .INIT(8'hb4)
  ) _240_ (
    .I0(Kgen),
    .I1(ki[54]),
    .I2(ki[22]),
    .O(_067_)
  );
LUT3  #(
    .INIT(8'hb4)
  ) _241_ (
    .I0(Kgen),
    .I1(ki[55]),
    .I2(ki[23]),
    .O(_068_)
  );
LUT4  #(
    .INIT(16'h8778)
  ) _242_ (
    .I0(ko[64]),
    .I1(Kgen),
    .I2(ki[0]),
    .I3(ki[32]),
    .O(ko[0])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _243_ (
    .I0(Kgen),
    .I1(so[0]),
    .I2(ki[64]),
    .I3(ki[96]),
    .O(ko[64])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _244_ (
    .I0(ko[65]),
    .I1(Kgen),
    .I2(ki[1]),
    .I3(ki[33]),
    .O(ko[1])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _245_ (
    .I0(Kgen),
    .I1(so[1]),
    .I2(ki[65]),
    .I3(ki[97]),
    .O(ko[65])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _246_ (
    .I0(ko[66]),
    .I1(Kgen),
    .I2(ki[2]),
    .I3(ki[34]),
    .O(ko[2])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _247_ (
    .I0(Kgen),
    .I1(so[2]),
    .I2(ki[66]),
    .I3(ki[98]),
    .O(ko[66])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _248_ (
    .I0(ko[67]),
    .I1(Kgen),
    .I2(ki[3]),
    .I3(ki[35]),
    .O(ko[3])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _249_ (
    .I0(Kgen),
    .I1(so[3]),
    .I2(ki[67]),
    .I3(ki[99]),
    .O(ko[67])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _250_ (
    .I0(ko[68]),
    .I1(Kgen),
    .I2(ki[4]),
    .I3(ki[36]),
    .O(ko[4])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _251_ (
    .I0(Kgen),
    .I1(so[4]),
    .I2(ki[68]),
    .I3(ki[100]),
    .O(ko[68])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _252_ (
    .I0(ko[69]),
    .I1(Kgen),
    .I2(ki[5]),
    .I3(ki[37]),
    .O(ko[5])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _253_ (
    .I0(Kgen),
    .I1(so[5]),
    .I2(ki[69]),
    .I3(ki[101]),
    .O(ko[69])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _254_ (
    .I0(ko[70]),
    .I1(Kgen),
    .I2(ki[6]),
    .I3(ki[38]),
    .O(ko[6])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _255_ (
    .I0(Kgen),
    .I1(so[6]),
    .I2(ki[70]),
    .I3(ki[102]),
    .O(ko[70])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _256_ (
    .I0(ko[71]),
    .I1(Kgen),
    .I2(ki[7]),
    .I3(ki[39]),
    .O(ko[7])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _257_ (
    .I0(Kgen),
    .I1(so[7]),
    .I2(ki[71]),
    .I3(ki[103]),
    .O(ko[71])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _258_ (
    .I0(ko[72]),
    .I1(Kgen),
    .I2(ki[8]),
    .I3(ki[40]),
    .O(ko[8])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _259_ (
    .I0(Kgen),
    .I1(so[8]),
    .I2(ki[72]),
    .I3(ki[104]),
    .O(ko[72])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _260_ (
    .I0(ko[73]),
    .I1(Kgen),
    .I2(ki[9]),
    .I3(ki[41]),
    .O(ko[9])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _261_ (
    .I0(Kgen),
    .I1(so[9]),
    .I2(ki[73]),
    .I3(ki[105]),
    .O(ko[73])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _262_ (
    .I0(ko[74]),
    .I1(Kgen),
    .I2(ki[10]),
    .I3(ki[42]),
    .O(ko[10])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _263_ (
    .I0(Kgen),
    .I1(so[10]),
    .I2(ki[74]),
    .I3(ki[106]),
    .O(ko[74])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _264_ (
    .I0(ko[75]),
    .I1(Kgen),
    .I2(ki[11]),
    .I3(ki[43]),
    .O(ko[11])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _265_ (
    .I0(Kgen),
    .I1(so[11]),
    .I2(ki[75]),
    .I3(ki[107]),
    .O(ko[75])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _266_ (
    .I0(ko[76]),
    .I1(Kgen),
    .I2(ki[12]),
    .I3(ki[44]),
    .O(ko[12])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _267_ (
    .I0(Kgen),
    .I1(so[12]),
    .I2(ki[76]),
    .I3(ki[108]),
    .O(ko[76])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _268_ (
    .I0(ko[77]),
    .I1(Kgen),
    .I2(ki[13]),
    .I3(ki[45]),
    .O(ko[13])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _269_ (
    .I0(Kgen),
    .I1(so[13]),
    .I2(ki[77]),
    .I3(ki[109]),
    .O(ko[77])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _270_ (
    .I0(ko[78]),
    .I1(Kgen),
    .I2(ki[14]),
    .I3(ki[46]),
    .O(ko[14])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _271_ (
    .I0(Kgen),
    .I1(so[14]),
    .I2(ki[78]),
    .I3(ki[110]),
    .O(ko[78])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _272_ (
    .I0(ko[79]),
    .I1(Kgen),
    .I2(ki[15]),
    .I3(ki[47]),
    .O(ko[15])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _273_ (
    .I0(Kgen),
    .I1(so[15]),
    .I2(ki[79]),
    .I3(ki[111]),
    .O(ko[79])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _274_ (
    .I0(ko[80]),
    .I1(Kgen),
    .I2(ki[16]),
    .I3(ki[48]),
    .O(ko[16])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _275_ (
    .I0(Kgen),
    .I1(so[16]),
    .I2(ki[80]),
    .I3(ki[112]),
    .O(ko[80])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _276_ (
    .I0(ko[81]),
    .I1(Kgen),
    .I2(ki[17]),
    .I3(ki[49]),
    .O(ko[17])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _277_ (
    .I0(Kgen),
    .I1(so[17]),
    .I2(ki[81]),
    .I3(ki[113]),
    .O(ko[81])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _278_ (
    .I0(ko[82]),
    .I1(Kgen),
    .I2(ki[18]),
    .I3(ki[50]),
    .O(ko[18])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _279_ (
    .I0(Kgen),
    .I1(so[18]),
    .I2(ki[82]),
    .I3(ki[114]),
    .O(ko[82])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _280_ (
    .I0(ko[83]),
    .I1(Kgen),
    .I2(ki[19]),
    .I3(ki[51]),
    .O(ko[19])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _281_ (
    .I0(Kgen),
    .I1(so[19]),
    .I2(ki[83]),
    .I3(ki[115]),
    .O(ko[83])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _282_ (
    .I0(ko[84]),
    .I1(Kgen),
    .I2(ki[20]),
    .I3(ki[52]),
    .O(ko[20])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _283_ (
    .I0(Kgen),
    .I1(so[20]),
    .I2(ki[84]),
    .I3(ki[116]),
    .O(ko[84])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _284_ (
    .I0(ko[85]),
    .I1(Kgen),
    .I2(ki[21]),
    .I3(ki[53]),
    .O(ko[21])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _285_ (
    .I0(Kgen),
    .I1(so[21]),
    .I2(ki[85]),
    .I3(ki[117]),
    .O(ko[85])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _286_ (
    .I0(ko[86]),
    .I1(Kgen),
    .I2(ki[22]),
    .I3(ki[54]),
    .O(ko[22])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _287_ (
    .I0(Kgen),
    .I1(so[22]),
    .I2(ki[86]),
    .I3(ki[118]),
    .O(ko[86])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _288_ (
    .I0(ko[87]),
    .I1(Kgen),
    .I2(ki[23]),
    .I3(ki[55]),
    .O(ko[23])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _289_ (
    .I0(Kgen),
    .I1(so[23]),
    .I2(ki[87]),
    .I3(ki[119]),
    .O(ko[87])
  );
LUT6  #(
    .INIT(64'h0f7fff8fff8f0f7f)
  ) _290_ (
    .I0(_000_[0]),
    .I1(Rrg[8]),
    .I2(Kgen),
    .I3(Rrg[0]),
    .I4(ki[88]),
    .I5(ki[120]),
    .O(_003_)
  );
LUT6  #(
    .INIT(64'hff8f0f7f0f7fff8f)
  ) _291_ (
    .I0(_000_[0]),
    .I1(Rrg[8]),
    .I2(Kgen),
    .I3(Rrg[0]),
    .I4(ki[88]),
    .I5(ki[120]),
    .O(_004_)
  );
MUXF7  _292_ (
    .I0(_003_),
    .I1(_004_),
    .O(_001_),
    .S(so[24])
  );
LUT6  #(
    .INIT(64'hf08000700070f080)
  ) _293_ (
    .I0(_000_[0]),
    .I1(Rrg[8]),
    .I2(Kgen),
    .I3(Rrg[0]),
    .I4(ki[88]),
    .I5(ki[120]),
    .O(_005_)
  );
LUT6  #(
    .INIT(64'h0070f080f0800070)
  ) _294_ (
    .I0(_000_[0]),
    .I1(Rrg[8]),
    .I2(Kgen),
    .I3(Rrg[0]),
    .I4(ki[88]),
    .I5(ki[120]),
    .O(_006_)
  );
MUXF7  _295_ (
    .I0(_005_),
    .I1(_006_),
    .O(_002_),
    .S(so[24])
  );
MUXF8  _296_ (
    .I0(_001_),
    .I1(_002_),
    .O(ko[24]),
    .S(_000_[7])
  );
LUT2  #(
    .INIT(4'h9)
  ) _297_ (
    .I0(ki[24]),
    .I1(ki[56]),
    .O(_000_[7])
  );
LUT6  #(
    .INIT(64'h0000000000000001)
  ) _298_ (
    .I0(Rrg[7]),
    .I1(Rrg[6]),
    .I2(Rrg[5]),
    .I3(Rrg[4]),
    .I4(Rrg[3]),
    .I5(Rrg[2]),
    .O(_007_)
  );
MUXF7  _299_ (
    .I0(_007_),
    .I1(1'h0),
    .O(_000_[0]),
    .S(Rrg[1])
  );
LUT6  #(
    .INIT(64'h28828228d77d7dd7)
  ) _300_ (
    .I0(Kgen),
    .I1(_078_[1]),
    .I2(ki[89]),
    .I3(ki[121]),
    .I4(so[25]),
    .I5(_081_[5]),
    .O(ko[25])
  );
LUT2  #(
    .INIT(4'h9)
  ) _301_ (
    .I0(ki[25]),
    .I1(ki[57]),
    .O(_081_[5])
  );
LUT6  #(
    .INIT(64'h0000000000000001)
  ) _302_ (
    .I0(Rrg[6]),
    .I1(Rrg[5]),
    .I2(Rrg[4]),
    .I3(Rrg[3]),
    .I4(Rrg[2]),
    .I5(Rrg[7]),
    .O(_010_)
  );
MUXF7  _303_ (
    .I0(_010_),
    .I1(1'h1),
    .O(_008_),
    .S(Rrg[1])
  );
MUXF7  _304_ (
    .I0(1'h0),
    .I1(1'h0),
    .O(_009_),
    .S(Rrg[1])
  );
MUXF8  _305_ (
    .I0(_008_),
    .I1(_009_),
    .O(_078_[1]),
    .S(Rrg[0])
  );
LUT6  #(
    .INIT(64'h75dfdf75df7575df)
  ) _306_ (
    .I0(Kgen),
    .I1(_011_[1]),
    .I2(_011_[2]),
    .I3(ki[90]),
    .I4(ki[122]),
    .I5(so[26]),
    .O(_012_)
  );
LUT6  #(
    .INIT(64'h8a20208a208a8a20)
  ) _307_ (
    .I0(Kgen),
    .I1(_011_[1]),
    .I2(_011_[2]),
    .I3(ki[90]),
    .I4(ki[122]),
    .I5(so[26]),
    .O(_013_)
  );
MUXF7  _308_ (
    .I0(_012_),
    .I1(_013_),
    .O(ko[26]),
    .S(_011_[6])
  );
LUT2  #(
    .INIT(4'h9)
  ) _309_ (
    .I0(ki[26]),
    .I1(ki[58]),
    .O(_011_[6])
  );
LUT6  #(
    .INIT(64'hfffffffffffffffe)
  ) _310_ (
    .I0(Rrg[7]),
    .I1(Rrg[6]),
    .I2(Rrg[5]),
    .I3(Rrg[4]),
    .I4(Rrg[3]),
    .I5(Rrg[8]),
    .O(_014_)
  );
MUXF7  _311_ (
    .I0(_014_),
    .I1(1'h0),
    .O(_011_[1]),
    .S(Rrg[2])
  );
LUT2  #(
    .INIT(4'h1)
  ) _312_ (
    .I0(Rrg[1]),
    .I1(Rrg[0]),
    .O(_011_[2])
  );
LUT6  #(
    .INIT(64'h75dfdf75df7575df)
  ) _313_ (
    .I0(Kgen),
    .I1(_015_[1]),
    .I2(_015_[2]),
    .I3(ki[91]),
    .I4(ki[123]),
    .I5(so[27]),
    .O(_016_)
  );
LUT6  #(
    .INIT(64'h8a20208a208a8a20)
  ) _314_ (
    .I0(Kgen),
    .I1(_015_[1]),
    .I2(_015_[2]),
    .I3(ki[91]),
    .I4(ki[123]),
    .I5(so[27]),
    .O(_017_)
  );
MUXF7  _315_ (
    .I0(_016_),
    .I1(_017_),
    .O(ko[27]),
    .S(_015_[6])
  );
LUT2  #(
    .INIT(4'h9)
  ) _316_ (
    .I0(ki[27]),
    .I1(ki[59]),
    .O(_015_[6])
  );
LUT6  #(
    .INIT(64'h00000000fffeffff)
  ) _317_ (
    .I0(Rrg[7]),
    .I1(Rrg[6]),
    .I2(Rrg[5]),
    .I3(Rrg[4]),
    .I4(Rrg[8]),
    .I5(Rrg[3]),
    .O(_015_[1])
  );
LUT3  #(
    .INIT(8'h01)
  ) _318_ (
    .I0(Rrg[2]),
    .I1(Rrg[1]),
    .I2(Rrg[0]),
    .O(_015_[2])
  );
LUT6  #(
    .INIT(64'h28828228d77d7dd7)
  ) _319_ (
    .I0(Kgen),
    .I1(_077_[1]),
    .I2(ki[92]),
    .I3(ki[124]),
    .I4(so[28]),
    .I5(_080_[5]),
    .O(ko[28])
  );
LUT2  #(
    .INIT(4'h9)
  ) _320_ (
    .I0(ki[28]),
    .I1(ki[60]),
    .O(_080_[5])
  );
LUT6  #(
    .INIT(64'h000000000000ff01)
  ) _321_ (
    .I0(Rrg[6]),
    .I1(Rrg[5]),
    .I2(Rrg[7]),
    .I3(Rrg[4]),
    .I4(Rrg[3]),
    .I5(Rrg[2]),
    .O(_020_)
  );
MUXF7  _322_ (
    .I0(_020_),
    .I1(1'h0),
    .O(_018_),
    .S(Rrg[1])
  );
MUXF7  _323_ (
    .I0(1'h0),
    .I1(1'h0),
    .O(_019_),
    .S(Rrg[1])
  );
MUXF8  _324_ (
    .I0(_018_),
    .I1(_019_),
    .O(_077_[1]),
    .S(Rrg[0])
  );
LUT6  #(
    .INIT(64'h75dfdf75df7575df)
  ) _325_ (
    .I0(Kgen),
    .I1(_021_[1]),
    .I2(_021_[2]),
    .I3(ki[93]),
    .I4(ki[125]),
    .I5(so[29]),
    .O(_022_)
  );
LUT6  #(
    .INIT(64'h8a20208a208a8a20)
  ) _326_ (
    .I0(Kgen),
    .I1(_021_[1]),
    .I2(_021_[2]),
    .I3(ki[93]),
    .I4(ki[125]),
    .I5(so[29]),
    .O(_023_)
  );
MUXF7  _327_ (
    .I0(_022_),
    .I1(_023_),
    .O(ko[29]),
    .S(_021_[6])
  );
LUT2  #(
    .INIT(4'h9)
  ) _328_ (
    .I0(ki[29]),
    .I1(ki[61]),
    .O(_021_[6])
  );
LUT4  #(
    .INIT(16'h00fe)
  ) _329_ (
    .I0(Rrg[7]),
    .I1(Rrg[6]),
    .I2(Rrg[8]),
    .I3(Rrg[5]),
    .O(_021_[1])
  );
LUT5  #(
    .INIT(32'd1)
  ) _330_ (
    .I0(Rrg[4]),
    .I1(Rrg[3]),
    .I2(Rrg[2]),
    .I3(Rrg[1]),
    .I4(Rrg[0]),
    .O(_021_[2])
  );
LUT6  #(
    .INIT(64'h28828228d77d7dd7)
  ) _331_ (
    .I0(Kgen),
    .I1(_076_[1]),
    .I2(ki[94]),
    .I3(ki[126]),
    .I4(so[30]),
    .I5(_079_[5]),
    .O(ko[30])
  );
LUT2  #(
    .INIT(4'h9)
  ) _332_ (
    .I0(ki[30]),
    .I1(ki[62]),
    .O(_079_[5])
  );
LUT6  #(
    .INIT(64'h0000000000000001)
  ) _333_ (
    .I0(Rrg[5]),
    .I1(Rrg[4]),
    .I2(Rrg[3]),
    .I3(Rrg[2]),
    .I4(Rrg[1]),
    .I5(Rrg[0]),
    .O(_024_)
  );
MUXF7  _334_ (
    .I0(1'h0),
    .I1(_024_),
    .O(_076_[1]),
    .S(Rrg[6])
  );
LUT6  #(
    .INIT(64'hd57f7fd57fd5d57f)
  ) _335_ (
    .I0(Kgen),
    .I1(_021_[2]),
    .I2(_025_[2]),
    .I3(ki[95]),
    .I4(ki[127]),
    .I5(so[31]),
    .O(_026_)
  );
LUT6  #(
    .INIT(64'h2a80802a802a2a80)
  ) _336_ (
    .I0(Kgen),
    .I1(_021_[2]),
    .I2(_025_[2]),
    .I3(ki[95]),
    .I4(ki[127]),
    .I5(so[31]),
    .O(_027_)
  );
MUXF7  _337_ (
    .I0(_026_),
    .I1(_027_),
    .O(ko[31]),
    .S(_025_[6])
  );
LUT2  #(
    .INIT(4'h9)
  ) _338_ (
    .I0(ki[31]),
    .I1(ki[63]),
    .O(_025_[6])
  );
LUT3  #(
    .INIT(8'h10)
  ) _339_ (
    .I0(Rrg[6]),
    .I1(Rrg[5]),
    .I2(Rrg[7]),
    .O(_025_[2])
  );
LUT6  #(
    .INIT(64'hff8f0f7f0070f080)
  ) _340_ (
    .I0(_000_[0]),
    .I1(Rrg[8]),
    .I2(Kgen),
    .I3(Rrg[0]),
    .I4(so[24]),
    .I5(ki[88]),
    .O(_028_)
  );
LUT6  #(
    .INIT(64'h0070f080ff8f0f7f)
  ) _341_ (
    .I0(_000_[0]),
    .I1(Rrg[8]),
    .I2(Kgen),
    .I3(Rrg[0]),
    .I4(so[24]),
    .I5(ki[88]),
    .O(_029_)
  );
MUXF7  _342_ (
    .I0(_028_),
    .I1(_029_),
    .O(ko[88]),
    .S(ki[120])
  );
LUT5  #(
    .INIT(32'd685233960)
  ) _343_ (
    .I0(Kgen),
    .I1(_078_[1]),
    .I2(so[25]),
    .I3(ki[89]),
    .I4(ki[121]),
    .O(ko[89])
  );
LUT6  #(
    .INIT(64'hb0404fbf4fbfb040)
  ) _344_ (
    .I0(_011_[1]),
    .I1(_011_[2]),
    .I2(Kgen),
    .I3(so[26]),
    .I4(ki[90]),
    .I5(ki[122]),
    .O(ko[90])
  );
LUT6  #(
    .INIT(64'hb0404fbf4fbfb040)
  ) _345_ (
    .I0(_015_[1]),
    .I1(_015_[2]),
    .I2(Kgen),
    .I3(so[27]),
    .I4(ki[91]),
    .I5(ki[123]),
    .O(ko[91])
  );
LUT5  #(
    .INIT(32'd685233960)
  ) _346_ (
    .I0(Kgen),
    .I1(_077_[1]),
    .I2(so[28]),
    .I3(ki[92]),
    .I4(ki[124]),
    .O(ko[92])
  );
LUT6  #(
    .INIT(64'hb0404fbf4fbfb040)
  ) _347_ (
    .I0(_021_[1]),
    .I1(_021_[2]),
    .I2(Kgen),
    .I3(so[29]),
    .I4(ki[93]),
    .I5(ki[125]),
    .O(ko[93])
  );
LUT5  #(
    .INIT(32'd685233960)
  ) _348_ (
    .I0(Kgen),
    .I1(_076_[1]),
    .I2(so[30]),
    .I3(ki[94]),
    .I4(ki[126]),
    .O(ko[94])
  );
LUT6  #(
    .INIT(64'h70808f7f8f7f7080)
  ) _349_ (
    .I0(_021_[2]),
    .I1(_025_[2]),
    .I2(Kgen),
    .I3(so[31]),
    .I4(ki[95]),
    .I5(ki[127]),
    .O(ko[95])
  );
LUT2  #(
    .INIT(4'h6)
  ) _350_ (
    .I0(ki[96]),
    .I1(so[0]),
    .O(ko[96])
  );
LUT2  #(
    .INIT(4'h6)
  ) _351_ (
    .I0(ki[97]),
    .I1(so[1]),
    .O(ko[97])
  );
LUT2  #(
    .INIT(4'h6)
  ) _352_ (
    .I0(ki[98]),
    .I1(so[2]),
    .O(ko[98])
  );
LUT2  #(
    .INIT(4'h6)
  ) _353_ (
    .I0(ki[99]),
    .I1(so[3]),
    .O(ko[99])
  );
LUT2  #(
    .INIT(4'h6)
  ) _354_ (
    .I0(ki[100]),
    .I1(so[4]),
    .O(ko[100])
  );
LUT2  #(
    .INIT(4'h6)
  ) _355_ (
    .I0(ki[101]),
    .I1(so[5]),
    .O(ko[101])
  );
LUT2  #(
    .INIT(4'h6)
  ) _356_ (
    .I0(ki[102]),
    .I1(so[6]),
    .O(ko[102])
  );
LUT2  #(
    .INIT(4'h6)
  ) _357_ (
    .I0(ki[103]),
    .I1(so[7]),
    .O(ko[103])
  );
LUT2  #(
    .INIT(4'h6)
  ) _358_ (
    .I0(ki[104]),
    .I1(so[8]),
    .O(ko[104])
  );
LUT2  #(
    .INIT(4'h6)
  ) _359_ (
    .I0(ki[105]),
    .I1(so[9]),
    .O(ko[105])
  );
LUT2  #(
    .INIT(4'h6)
  ) _360_ (
    .I0(ki[106]),
    .I1(so[10]),
    .O(ko[106])
  );
LUT2  #(
    .INIT(4'h6)
  ) _361_ (
    .I0(ki[107]),
    .I1(so[11]),
    .O(ko[107])
  );
LUT2  #(
    .INIT(4'h6)
  ) _362_ (
    .I0(ki[108]),
    .I1(so[12]),
    .O(ko[108])
  );
LUT2  #(
    .INIT(4'h6)
  ) _363_ (
    .I0(ki[109]),
    .I1(so[13]),
    .O(ko[109])
  );
LUT2  #(
    .INIT(4'h6)
  ) _364_ (
    .I0(ki[110]),
    .I1(so[14]),
    .O(ko[110])
  );
LUT2  #(
    .INIT(4'h6)
  ) _365_ (
    .I0(ki[111]),
    .I1(so[15]),
    .O(ko[111])
  );
LUT2  #(
    .INIT(4'h6)
  ) _366_ (
    .I0(ki[112]),
    .I1(so[16]),
    .O(ko[112])
  );
LUT2  #(
    .INIT(4'h6)
  ) _367_ (
    .I0(ki[113]),
    .I1(so[17]),
    .O(ko[113])
  );
LUT2  #(
    .INIT(4'h6)
  ) _368_ (
    .I0(ki[114]),
    .I1(so[18]),
    .O(ko[114])
  );
LUT2  #(
    .INIT(4'h6)
  ) _369_ (
    .I0(ki[115]),
    .I1(so[19]),
    .O(ko[115])
  );
LUT2  #(
    .INIT(4'h6)
  ) _370_ (
    .I0(ki[116]),
    .I1(so[20]),
    .O(ko[116])
  );
LUT2  #(
    .INIT(4'h6)
  ) _371_ (
    .I0(ki[117]),
    .I1(so[21]),
    .O(ko[117])
  );
LUT2  #(
    .INIT(4'h6)
  ) _372_ (
    .I0(ki[118]),
    .I1(so[22]),
    .O(ko[118])
  );
LUT2  #(
    .INIT(4'h6)
  ) _373_ (
    .I0(ki[119]),
    .I1(so[23]),
    .O(ko[119])
  );
LUT5  #(
    .INIT(32'd4161210360)
  ) _374_ (
    .I0(_000_[0]),
    .I1(Rrg[8]),
    .I2(Rrg[0]),
    .I3(ki[120]),
    .I4(so[24]),
    .O(ko[120])
  );
LUT3  #(
    .INIT(8'h96)
  ) _375_ (
    .I0(_078_[1]),
    .I1(ki[121]),
    .I2(so[25]),
    .O(ko[121])
  );
LUT4  #(
    .INIT(16'h4bb4)
  ) _376_ (
    .I0(_011_[1]),
    .I1(_011_[2]),
    .I2(ki[122]),
    .I3(so[26]),
    .O(ko[122])
  );
LUT4  #(
    .INIT(16'h4bb4)
  ) _377_ (
    .I0(_015_[1]),
    .I1(_015_[2]),
    .I2(ki[123]),
    .I3(so[27]),
    .O(ko[123])
  );
LUT3  #(
    .INIT(8'h96)
  ) _378_ (
    .I0(_077_[1]),
    .I1(ki[124]),
    .I2(so[28]),
    .O(ko[124])
  );
LUT4  #(
    .INIT(16'h4bb4)
  ) _379_ (
    .I0(_021_[1]),
    .I1(_021_[2]),
    .I2(ki[125]),
    .I3(so[29]),
    .O(ko[125])
  );
LUT3  #(
    .INIT(8'h96)
  ) _380_ (
    .I0(_076_[1]),
    .I1(ki[126]),
    .I2(so[30]),
    .O(ko[126])
  );
LUT4  #(
    .INIT(16'h8778)
  ) _381_ (
    .I0(_021_[2]),
    .I1(_025_[2]),
    .I2(ki[127]),
    .I3(so[31]),
    .O(ko[127])
  );
LUT2  #(
    .INIT(4'h6)
  ) _382_ (
    .I0(ki[0]),
    .I1(sb[0]),
    .O(\do [0])
  );
LUT2  #(
    .INIT(4'h6)
  ) _383_ (
    .I0(ki[1]),
    .I1(sb[1]),
    .O(\do [1])
  );
LUT2  #(
    .INIT(4'h6)
  ) _384_ (
    .I0(ki[2]),
    .I1(sb[2]),
    .O(\do [2])
  );
LUT2  #(
    .INIT(4'h6)
  ) _385_ (
    .I0(ki[3]),
    .I1(sb[3]),
    .O(\do [3])
  );
LUT2  #(
    .INIT(4'h6)
  ) _386_ (
    .I0(ki[4]),
    .I1(sb[4]),
    .O(\do [4])
  );
LUT2  #(
    .INIT(4'h6)
  ) _387_ (
    .I0(ki[5]),
    .I1(sb[5]),
    .O(\do [5])
  );
LUT2  #(
    .INIT(4'h6)
  ) _388_ (
    .I0(ki[6]),
    .I1(sb[6]),
    .O(\do [6])
  );
LUT2  #(
    .INIT(4'h6)
  ) _389_ (
    .I0(ki[7]),
    .I1(sb[7]),
    .O(\do [7])
  );
LUT2  #(
    .INIT(4'h6)
  ) _390_ (
    .I0(ki[8]),
    .I1(sb[8]),
    .O(\do [8])
  );
LUT2  #(
    .INIT(4'h6)
  ) _391_ (
    .I0(ki[9]),
    .I1(sb[9]),
    .O(\do [9])
  );
LUT2  #(
    .INIT(4'h6)
  ) _392_ (
    .I0(ki[10]),
    .I1(sb[10]),
    .O(\do [10])
  );
LUT2  #(
    .INIT(4'h6)
  ) _393_ (
    .I0(ki[11]),
    .I1(sb[11]),
    .O(\do [11])
  );
LUT2  #(
    .INIT(4'h6)
  ) _394_ (
    .I0(ki[12]),
    .I1(sb[12]),
    .O(\do [12])
  );
LUT2  #(
    .INIT(4'h6)
  ) _395_ (
    .I0(ki[13]),
    .I1(sb[13]),
    .O(\do [13])
  );
LUT2  #(
    .INIT(4'h6)
  ) _396_ (
    .I0(ki[14]),
    .I1(sb[14]),
    .O(\do [14])
  );
LUT2  #(
    .INIT(4'h6)
  ) _397_ (
    .I0(ki[15]),
    .I1(sb[15]),
    .O(\do [15])
  );
LUT2  #(
    .INIT(4'h6)
  ) _398_ (
    .I0(ki[16]),
    .I1(sb[16]),
    .O(\do [16])
  );
LUT2  #(
    .INIT(4'h6)
  ) _399_ (
    .I0(ki[17]),
    .I1(sb[17]),
    .O(\do [17])
  );
LUT2  #(
    .INIT(4'h6)
  ) _400_ (
    .I0(ki[18]),
    .I1(sb[18]),
    .O(\do [18])
  );
LUT2  #(
    .INIT(4'h6)
  ) _401_ (
    .I0(ki[19]),
    .I1(sb[19]),
    .O(\do [19])
  );
LUT2  #(
    .INIT(4'h6)
  ) _402_ (
    .I0(ki[20]),
    .I1(sb[20]),
    .O(\do [20])
  );
LUT2  #(
    .INIT(4'h6)
  ) _403_ (
    .I0(ki[21]),
    .I1(sb[21]),
    .O(\do [21])
  );
LUT2  #(
    .INIT(4'h6)
  ) _404_ (
    .I0(ki[22]),
    .I1(sb[22]),
    .O(\do [22])
  );
LUT2  #(
    .INIT(4'h6)
  ) _405_ (
    .I0(ki[23]),
    .I1(sb[23]),
    .O(\do [23])
  );
LUT2  #(
    .INIT(4'h6)
  ) _406_ (
    .I0(ki[24]),
    .I1(sb[24]),
    .O(\do [24])
  );
LUT2  #(
    .INIT(4'h6)
  ) _407_ (
    .I0(ki[25]),
    .I1(sb[25]),
    .O(\do [25])
  );
LUT2  #(
    .INIT(4'h6)
  ) _408_ (
    .I0(ki[26]),
    .I1(sb[26]),
    .O(\do [26])
  );
LUT2  #(
    .INIT(4'h6)
  ) _409_ (
    .I0(ki[27]),
    .I1(sb[27]),
    .O(\do [27])
  );
LUT2  #(
    .INIT(4'h6)
  ) _410_ (
    .I0(ki[28]),
    .I1(sb[28]),
    .O(\do [28])
  );
LUT2  #(
    .INIT(4'h6)
  ) _411_ (
    .I0(ki[29]),
    .I1(sb[29]),
    .O(\do [29])
  );
LUT2  #(
    .INIT(4'h6)
  ) _412_ (
    .I0(ki[30]),
    .I1(sb[30]),
    .O(\do [30])
  );
LUT2  #(
    .INIT(4'h6)
  ) _413_ (
    .I0(ki[31]),
    .I1(sb[31]),
    .O(\do [31])
  );
LUT2  #(
    .INIT(4'h6)
  ) _414_ (
    .I0(ki[32]),
    .I1(sb[32]),
    .O(\do [32])
  );
LUT2  #(
    .INIT(4'h6)
  ) _415_ (
    .I0(ki[33]),
    .I1(sb[33]),
    .O(\do [33])
  );
LUT2  #(
    .INIT(4'h6)
  ) _416_ (
    .I0(ki[34]),
    .I1(sb[34]),
    .O(\do [34])
  );
LUT2  #(
    .INIT(4'h6)
  ) _417_ (
    .I0(ki[35]),
    .I1(sb[35]),
    .O(\do [35])
  );
LUT2  #(
    .INIT(4'h6)
  ) _418_ (
    .I0(ki[36]),
    .I1(sb[36]),
    .O(\do [36])
  );
LUT2  #(
    .INIT(4'h6)
  ) _419_ (
    .I0(ki[37]),
    .I1(sb[37]),
    .O(\do [37])
  );
LUT2  #(
    .INIT(4'h6)
  ) _420_ (
    .I0(ki[38]),
    .I1(sb[38]),
    .O(\do [38])
  );
LUT2  #(
    .INIT(4'h6)
  ) _421_ (
    .I0(ki[39]),
    .I1(sb[39]),
    .O(\do [39])
  );
LUT2  #(
    .INIT(4'h6)
  ) _422_ (
    .I0(ki[40]),
    .I1(sb[40]),
    .O(\do [40])
  );
LUT2  #(
    .INIT(4'h6)
  ) _423_ (
    .I0(ki[41]),
    .I1(sb[41]),
    .O(\do [41])
  );
LUT2  #(
    .INIT(4'h6)
  ) _424_ (
    .I0(ki[42]),
    .I1(sb[42]),
    .O(\do [42])
  );
LUT2  #(
    .INIT(4'h6)
  ) _425_ (
    .I0(ki[43]),
    .I1(sb[43]),
    .O(\do [43])
  );
LUT2  #(
    .INIT(4'h6)
  ) _426_ (
    .I0(ki[44]),
    .I1(sb[44]),
    .O(\do [44])
  );
LUT2  #(
    .INIT(4'h6)
  ) _427_ (
    .I0(ki[45]),
    .I1(sb[45]),
    .O(\do [45])
  );
LUT2  #(
    .INIT(4'h6)
  ) _428_ (
    .I0(ki[46]),
    .I1(sb[46]),
    .O(\do [46])
  );
LUT2  #(
    .INIT(4'h6)
  ) _429_ (
    .I0(ki[47]),
    .I1(sb[47]),
    .O(\do [47])
  );
LUT2  #(
    .INIT(4'h6)
  ) _430_ (
    .I0(ki[48]),
    .I1(sb[48]),
    .O(\do [48])
  );
LUT2  #(
    .INIT(4'h6)
  ) _431_ (
    .I0(ki[49]),
    .I1(sb[49]),
    .O(\do [49])
  );
LUT2  #(
    .INIT(4'h6)
  ) _432_ (
    .I0(ki[50]),
    .I1(sb[50]),
    .O(\do [50])
  );
LUT2  #(
    .INIT(4'h6)
  ) _433_ (
    .I0(ki[51]),
    .I1(sb[51]),
    .O(\do [51])
  );
LUT2  #(
    .INIT(4'h6)
  ) _434_ (
    .I0(ki[52]),
    .I1(sb[52]),
    .O(\do [52])
  );
LUT2  #(
    .INIT(4'h6)
  ) _435_ (
    .I0(ki[53]),
    .I1(sb[53]),
    .O(\do [53])
  );
LUT2  #(
    .INIT(4'h6)
  ) _436_ (
    .I0(ki[54]),
    .I1(sb[54]),
    .O(\do [54])
  );
LUT2  #(
    .INIT(4'h6)
  ) _437_ (
    .I0(ki[55]),
    .I1(sb[55]),
    .O(\do [55])
  );
LUT2  #(
    .INIT(4'h6)
  ) _438_ (
    .I0(ki[56]),
    .I1(sb[56]),
    .O(\do [56])
  );
LUT2  #(
    .INIT(4'h6)
  ) _439_ (
    .I0(ki[57]),
    .I1(sb[57]),
    .O(\do [57])
  );
LUT2  #(
    .INIT(4'h6)
  ) _440_ (
    .I0(ki[58]),
    .I1(sb[58]),
    .O(\do [58])
  );
LUT2  #(
    .INIT(4'h6)
  ) _441_ (
    .I0(ki[59]),
    .I1(sb[59]),
    .O(\do [59])
  );
LUT2  #(
    .INIT(4'h6)
  ) _442_ (
    .I0(ki[60]),
    .I1(sb[60]),
    .O(\do [60])
  );
LUT2  #(
    .INIT(4'h6)
  ) _443_ (
    .I0(ki[61]),
    .I1(sb[61]),
    .O(\do [61])
  );
LUT2  #(
    .INIT(4'h6)
  ) _444_ (
    .I0(ki[62]),
    .I1(sb[62]),
    .O(\do [62])
  );
LUT2  #(
    .INIT(4'h6)
  ) _445_ (
    .I0(ki[63]),
    .I1(sb[63]),
    .O(\do [63])
  );
LUT2  #(
    .INIT(4'h6)
  ) _446_ (
    .I0(ki[64]),
    .I1(sb[64]),
    .O(\do [64])
  );
LUT2  #(
    .INIT(4'h6)
  ) _447_ (
    .I0(ki[65]),
    .I1(sb[65]),
    .O(\do [65])
  );
LUT2  #(
    .INIT(4'h6)
  ) _448_ (
    .I0(ki[66]),
    .I1(sb[66]),
    .O(\do [66])
  );
LUT2  #(
    .INIT(4'h6)
  ) _449_ (
    .I0(ki[67]),
    .I1(sb[67]),
    .O(\do [67])
  );
LUT2  #(
    .INIT(4'h6)
  ) _450_ (
    .I0(ki[68]),
    .I1(sb[68]),
    .O(\do [68])
  );
LUT2  #(
    .INIT(4'h6)
  ) _451_ (
    .I0(ki[69]),
    .I1(sb[69]),
    .O(\do [69])
  );
LUT2  #(
    .INIT(4'h6)
  ) _452_ (
    .I0(ki[70]),
    .I1(sb[70]),
    .O(\do [70])
  );
LUT2  #(
    .INIT(4'h6)
  ) _453_ (
    .I0(ki[71]),
    .I1(sb[71]),
    .O(\do [71])
  );
LUT2  #(
    .INIT(4'h6)
  ) _454_ (
    .I0(ki[72]),
    .I1(sb[72]),
    .O(\do [72])
  );
LUT2  #(
    .INIT(4'h6)
  ) _455_ (
    .I0(ki[73]),
    .I1(sb[73]),
    .O(\do [73])
  );
LUT2  #(
    .INIT(4'h6)
  ) _456_ (
    .I0(ki[74]),
    .I1(sb[74]),
    .O(\do [74])
  );
LUT2  #(
    .INIT(4'h6)
  ) _457_ (
    .I0(ki[75]),
    .I1(sb[75]),
    .O(\do [75])
  );
LUT2  #(
    .INIT(4'h6)
  ) _458_ (
    .I0(ki[76]),
    .I1(sb[76]),
    .O(\do [76])
  );
LUT2  #(
    .INIT(4'h6)
  ) _459_ (
    .I0(ki[77]),
    .I1(sb[77]),
    .O(\do [77])
  );
LUT2  #(
    .INIT(4'h6)
  ) _460_ (
    .I0(ki[78]),
    .I1(sb[78]),
    .O(\do [78])
  );
LUT2  #(
    .INIT(4'h6)
  ) _461_ (
    .I0(ki[79]),
    .I1(sb[79]),
    .O(\do [79])
  );
LUT2  #(
    .INIT(4'h6)
  ) _462_ (
    .I0(ki[80]),
    .I1(sb[80]),
    .O(\do [80])
  );
LUT2  #(
    .INIT(4'h6)
  ) _463_ (
    .I0(ki[81]),
    .I1(sb[81]),
    .O(\do [81])
  );
LUT2  #(
    .INIT(4'h6)
  ) _464_ (
    .I0(ki[82]),
    .I1(sb[82]),
    .O(\do [82])
  );
LUT2  #(
    .INIT(4'h6)
  ) _465_ (
    .I0(ki[83]),
    .I1(sb[83]),
    .O(\do [83])
  );
LUT2  #(
    .INIT(4'h6)
  ) _466_ (
    .I0(ki[84]),
    .I1(sb[84]),
    .O(\do [84])
  );
LUT2  #(
    .INIT(4'h6)
  ) _467_ (
    .I0(ki[85]),
    .I1(sb[85]),
    .O(\do [85])
  );
LUT2  #(
    .INIT(4'h6)
  ) _468_ (
    .I0(ki[86]),
    .I1(sb[86]),
    .O(\do [86])
  );
LUT2  #(
    .INIT(4'h6)
  ) _469_ (
    .I0(ki[87]),
    .I1(sb[87]),
    .O(\do [87])
  );
LUT2  #(
    .INIT(4'h6)
  ) _470_ (
    .I0(ki[88]),
    .I1(sb[88]),
    .O(\do [88])
  );
LUT2  #(
    .INIT(4'h6)
  ) _471_ (
    .I0(ki[89]),
    .I1(sb[89]),
    .O(\do [89])
  );
LUT2  #(
    .INIT(4'h6)
  ) _472_ (
    .I0(ki[90]),
    .I1(sb[90]),
    .O(\do [90])
  );
LUT2  #(
    .INIT(4'h6)
  ) _473_ (
    .I0(ki[91]),
    .I1(sb[91]),
    .O(\do [91])
  );
LUT2  #(
    .INIT(4'h6)
  ) _474_ (
    .I0(ki[92]),
    .I1(sb[92]),
    .O(\do [92])
  );
LUT2  #(
    .INIT(4'h6)
  ) _475_ (
    .I0(ki[93]),
    .I1(sb[93]),
    .O(\do [93])
  );
LUT2  #(
    .INIT(4'h6)
  ) _476_ (
    .I0(ki[94]),
    .I1(sb[94]),
    .O(\do [94])
  );
LUT2  #(
    .INIT(4'h6)
  ) _477_ (
    .I0(ki[95]),
    .I1(sb[95]),
    .O(\do [95])
  );
LUT2  #(
    .INIT(4'h6)
  ) _478_ (
    .I0(ki[96]),
    .I1(sb[96]),
    .O(\do [96])
  );
LUT2  #(
    .INIT(4'h6)
  ) _479_ (
    .I0(ki[97]),
    .I1(sb[97]),
    .O(\do [97])
  );
LUT2  #(
    .INIT(4'h6)
  ) _480_ (
    .I0(ki[98]),
    .I1(sb[98]),
    .O(\do [98])
  );
LUT2  #(
    .INIT(4'h6)
  ) _481_ (
    .I0(ki[99]),
    .I1(sb[99]),
    .O(\do [99])
  );
LUT2  #(
    .INIT(4'h6)
  ) _482_ (
    .I0(ki[100]),
    .I1(sb[100]),
    .O(\do [100])
  );
LUT2  #(
    .INIT(4'h6)
  ) _483_ (
    .I0(ki[101]),
    .I1(sb[101]),
    .O(\do [101])
  );
LUT2  #(
    .INIT(4'h6)
  ) _484_ (
    .I0(ki[102]),
    .I1(sb[102]),
    .O(\do [102])
  );
LUT2  #(
    .INIT(4'h6)
  ) _485_ (
    .I0(ki[103]),
    .I1(sb[103]),
    .O(\do [103])
  );
LUT2  #(
    .INIT(4'h6)
  ) _486_ (
    .I0(ki[104]),
    .I1(sb[104]),
    .O(\do [104])
  );
LUT2  #(
    .INIT(4'h6)
  ) _487_ (
    .I0(ki[105]),
    .I1(sb[105]),
    .O(\do [105])
  );
LUT2  #(
    .INIT(4'h6)
  ) _488_ (
    .I0(ki[106]),
    .I1(sb[106]),
    .O(\do [106])
  );
LUT2  #(
    .INIT(4'h6)
  ) _489_ (
    .I0(ki[107]),
    .I1(sb[107]),
    .O(\do [107])
  );
LUT2  #(
    .INIT(4'h6)
  ) _490_ (
    .I0(ki[108]),
    .I1(sb[108]),
    .O(\do [108])
  );
LUT2  #(
    .INIT(4'h6)
  ) _491_ (
    .I0(ki[109]),
    .I1(sb[109]),
    .O(\do [109])
  );
LUT2  #(
    .INIT(4'h6)
  ) _492_ (
    .I0(ki[110]),
    .I1(sb[110]),
    .O(\do [110])
  );
LUT2  #(
    .INIT(4'h6)
  ) _493_ (
    .I0(ki[111]),
    .I1(sb[111]),
    .O(\do [111])
  );
LUT2  #(
    .INIT(4'h6)
  ) _494_ (
    .I0(ki[112]),
    .I1(sb[112]),
    .O(\do [112])
  );
LUT2  #(
    .INIT(4'h6)
  ) _495_ (
    .I0(ki[113]),
    .I1(sb[113]),
    .O(\do [113])
  );
LUT2  #(
    .INIT(4'h6)
  ) _496_ (
    .I0(ki[114]),
    .I1(sb[114]),
    .O(\do [114])
  );
LUT2  #(
    .INIT(4'h6)
  ) _497_ (
    .I0(ki[115]),
    .I1(sb[115]),
    .O(\do [115])
  );
LUT2  #(
    .INIT(4'h6)
  ) _498_ (
    .I0(ki[116]),
    .I1(sb[116]),
    .O(\do [116])
  );
LUT2  #(
    .INIT(4'h6)
  ) _499_ (
    .I0(ki[117]),
    .I1(sb[117]),
    .O(\do [117])
  );
LUT2  #(
    .INIT(4'h6)
  ) _500_ (
    .I0(ki[118]),
    .I1(sb[118]),
    .O(\do [118])
  );
LUT2  #(
    .INIT(4'h6)
  ) _501_ (
    .I0(ki[119]),
    .I1(sb[119]),
    .O(\do [119])
  );
LUT2  #(
    .INIT(4'h6)
  ) _502_ (
    .I0(ki[120]),
    .I1(sb[120]),
    .O(\do [120])
  );
LUT2  #(
    .INIT(4'h6)
  ) _503_ (
    .I0(ki[121]),
    .I1(sb[121]),
    .O(\do [121])
  );
LUT2  #(
    .INIT(4'h6)
  ) _504_ (
    .I0(ki[122]),
    .I1(sb[122]),
    .O(\do [122])
  );
LUT2  #(
    .INIT(4'h6)
  ) _505_ (
    .I0(ki[123]),
    .I1(sb[123]),
    .O(\do [123])
  );
LUT2  #(
    .INIT(4'h6)
  ) _506_ (
    .I0(ki[124]),
    .I1(sb[124]),
    .O(\do [124])
  );
LUT2  #(
    .INIT(4'h6)
  ) _507_ (
    .I0(ki[125]),
    .I1(sb[125]),
    .O(\do [125])
  );
LUT2  #(
    .INIT(4'h6)
  ) _508_ (
    .I0(ki[126]),
    .I1(sb[126]),
    .O(\do [126])
  );
LUT2  #(
    .INIT(4'h6)
  ) _509_ (
    .I0(ki[127]),
    .I1(sb[127]),
    .O(\do [127])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _510_ (
    .I0(ko[64]),
    .I1(ki[64]),
    .I2(Kgen),
    .I3(ki[32]),
    .O(ko[32])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _511_ (
    .I0(ko[65]),
    .I1(ki[65]),
    .I2(Kgen),
    .I3(ki[33]),
    .O(ko[33])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _512_ (
    .I0(ko[66]),
    .I1(ki[66]),
    .I2(Kgen),
    .I3(ki[34]),
    .O(ko[34])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _513_ (
    .I0(ko[67]),
    .I1(ki[67]),
    .I2(Kgen),
    .I3(ki[35]),
    .O(ko[35])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _514_ (
    .I0(ko[68]),
    .I1(ki[68]),
    .I2(Kgen),
    .I3(ki[36]),
    .O(ko[36])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _515_ (
    .I0(ko[69]),
    .I1(ki[69]),
    .I2(Kgen),
    .I3(ki[37]),
    .O(ko[37])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _516_ (
    .I0(ko[70]),
    .I1(ki[70]),
    .I2(Kgen),
    .I3(ki[38]),
    .O(ko[38])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _517_ (
    .I0(ko[71]),
    .I1(ki[71]),
    .I2(Kgen),
    .I3(ki[39]),
    .O(ko[39])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _518_ (
    .I0(ko[72]),
    .I1(ki[72]),
    .I2(Kgen),
    .I3(ki[40]),
    .O(ko[40])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _519_ (
    .I0(ko[73]),
    .I1(ki[73]),
    .I2(Kgen),
    .I3(ki[41]),
    .O(ko[41])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _520_ (
    .I0(ko[74]),
    .I1(ki[74]),
    .I2(Kgen),
    .I3(ki[42]),
    .O(ko[42])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _521_ (
    .I0(ko[75]),
    .I1(ki[75]),
    .I2(Kgen),
    .I3(ki[43]),
    .O(ko[43])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _522_ (
    .I0(ko[76]),
    .I1(ki[76]),
    .I2(Kgen),
    .I3(ki[44]),
    .O(ko[44])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _523_ (
    .I0(ko[77]),
    .I1(ki[77]),
    .I2(Kgen),
    .I3(ki[45]),
    .O(ko[45])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _524_ (
    .I0(ko[78]),
    .I1(ki[78]),
    .I2(Kgen),
    .I3(ki[46]),
    .O(ko[46])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _525_ (
    .I0(ko[79]),
    .I1(ki[79]),
    .I2(Kgen),
    .I3(ki[47]),
    .O(ko[47])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _526_ (
    .I0(ko[80]),
    .I1(ki[80]),
    .I2(Kgen),
    .I3(ki[48]),
    .O(ko[48])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _527_ (
    .I0(ko[81]),
    .I1(ki[81]),
    .I2(Kgen),
    .I3(ki[49]),
    .O(ko[49])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _528_ (
    .I0(ko[82]),
    .I1(ki[82]),
    .I2(Kgen),
    .I3(ki[50]),
    .O(ko[50])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _529_ (
    .I0(ko[83]),
    .I1(ki[83]),
    .I2(Kgen),
    .I3(ki[51]),
    .O(ko[51])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _530_ (
    .I0(ko[84]),
    .I1(ki[84]),
    .I2(Kgen),
    .I3(ki[52]),
    .O(ko[52])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _531_ (
    .I0(ko[85]),
    .I1(ki[85]),
    .I2(Kgen),
    .I3(ki[53]),
    .O(ko[53])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _532_ (
    .I0(ko[86]),
    .I1(ki[86]),
    .I2(Kgen),
    .I3(ki[54]),
    .O(ko[54])
  );
LUT4  #(
    .INIT(16'h53ac)
  ) _533_ (
    .I0(ko[87]),
    .I1(ki[87]),
    .I2(Kgen),
    .I3(ki[55]),
    .O(ko[55])
  );
LUT6  #(
    .INIT(64'hf08000700070f080)
  ) _534_ (
    .I0(_000_[0]),
    .I1(Rrg[8]),
    .I2(Kgen),
    .I3(Rrg[0]),
    .I4(ki[120]),
    .I5(so[24]),
    .O(_032_)
  );
LUT6  #(
    .INIT(64'h0f7fff8fff8f0f7f)
  ) _535_ (
    .I0(_000_[0]),
    .I1(Rrg[8]),
    .I2(Kgen),
    .I3(Rrg[0]),
    .I4(ki[120]),
    .I5(so[24]),
    .O(_033_)
  );
MUXF7  _536_ (
    .I0(_032_),
    .I1(_033_),
    .O(_030_),
    .S(ki[88])
  );
LUT6  #(
    .INIT(64'h0f7fff8fff8f0f7f)
  ) _537_ (
    .I0(_000_[0]),
    .I1(Rrg[8]),
    .I2(Kgen),
    .I3(Rrg[0]),
    .I4(ki[120]),
    .I5(so[24]),
    .O(_034_)
  );
LUT6  #(
    .INIT(64'hf08000700070f080)
  ) _538_ (
    .I0(_000_[0]),
    .I1(Rrg[8]),
    .I2(Kgen),
    .I3(Rrg[0]),
    .I4(ki[120]),
    .I5(so[24]),
    .O(_035_)
  );
MUXF7  _539_ (
    .I0(_034_),
    .I1(_035_),
    .O(_031_),
    .S(ki[88])
  );
MUXF8  _540_ (
    .I0(_030_),
    .I1(_031_),
    .O(ko[56]),
    .S(ki[56])
  );
LUT6  #(
    .INIT(64'h82287dd77dd78228)
  ) _541_ (
    .I0(Kgen),
    .I1(_078_[1]),
    .I2(ki[121]),
    .I3(so[25]),
    .I4(ki[89]),
    .I5(ki[57]),
    .O(ko[57])
  );
LUT6  #(
    .INIT(64'hdf7575df208a8a20)
  ) _542_ (
    .I0(Kgen),
    .I1(_011_[1]),
    .I2(_011_[2]),
    .I3(ki[122]),
    .I4(so[26]),
    .I5(ki[90]),
    .O(_036_)
  );
LUT6  #(
    .INIT(64'h208a8a20df7575df)
  ) _543_ (
    .I0(Kgen),
    .I1(_011_[1]),
    .I2(_011_[2]),
    .I3(ki[122]),
    .I4(so[26]),
    .I5(ki[90]),
    .O(_037_)
  );
MUXF7  _544_ (
    .I0(_036_),
    .I1(_037_),
    .O(ko[58]),
    .S(ki[58])
  );
LUT6  #(
    .INIT(64'hdf7575df208a8a20)
  ) _545_ (
    .I0(Kgen),
    .I1(_015_[1]),
    .I2(_015_[2]),
    .I3(ki[123]),
    .I4(so[27]),
    .I5(ki[91]),
    .O(_038_)
  );
LUT6  #(
    .INIT(64'h208a8a20df7575df)
  ) _546_ (
    .I0(Kgen),
    .I1(_015_[1]),
    .I2(_015_[2]),
    .I3(ki[123]),
    .I4(so[27]),
    .I5(ki[91]),
    .O(_039_)
  );
MUXF7  _547_ (
    .I0(_038_),
    .I1(_039_),
    .O(ko[59]),
    .S(ki[59])
  );
LUT6  #(
    .INIT(64'h82287dd77dd78228)
  ) _548_ (
    .I0(Kgen),
    .I1(_077_[1]),
    .I2(ki[124]),
    .I3(so[28]),
    .I4(ki[92]),
    .I5(ki[60]),
    .O(ko[60])
  );
LUT6  #(
    .INIT(64'hdf7575df208a8a20)
  ) _549_ (
    .I0(Kgen),
    .I1(_021_[1]),
    .I2(_021_[2]),
    .I3(ki[125]),
    .I4(so[29]),
    .I5(ki[93]),
    .O(_040_)
  );
LUT6  #(
    .INIT(64'h208a8a20df7575df)
  ) _550_ (
    .I0(Kgen),
    .I1(_021_[1]),
    .I2(_021_[2]),
    .I3(ki[125]),
    .I4(so[29]),
    .I5(ki[93]),
    .O(_041_)
  );
MUXF7  _551_ (
    .I0(_040_),
    .I1(_041_),
    .O(ko[61]),
    .S(ki[61])
  );
LUT6  #(
    .INIT(64'h82287dd77dd78228)
  ) _552_ (
    .I0(Kgen),
    .I1(_076_[1]),
    .I2(ki[126]),
    .I3(so[30]),
    .I4(ki[94]),
    .I5(ki[62]),
    .O(ko[62])
  );
LUT6  #(
    .INIT(64'h7fd5d57f802a2a80)
  ) _553_ (
    .I0(Kgen),
    .I1(_021_[2]),
    .I2(_025_[2]),
    .I3(ki[127]),
    .I4(so[31]),
    .I5(ki[95]),
    .O(_042_)
  );
LUT6  #(
    .INIT(64'h802a2a807fd5d57f)
  ) _554_ (
    .I0(Kgen),
    .I1(_021_[2]),
    .I2(_025_[2]),
    .I3(ki[127]),
    .I4(so[31]),
    .I5(ki[95]),
    .O(_043_)
  );
MUXF7  _555_ (
    .I0(_042_),
    .I1(_043_),
    .O(ko[63]),
    .S(ki[63])
  );
AES_Comp_InvMixColumns  MX0 (
    .x(di[31:0]),
    .y(mx[31:0])
  );
AES_Comp_InvMixColumns  MX1 (
    .x(di[63:32]),
    .y(mx[63:32])
  );
AES_Comp_InvMixColumns  MX2 (
    .x(di[95:64]),
    .y(mx[95:64])
  );
AES_Comp_InvMixColumns  MX3 (
    .x(di[127:96]),
    .y(mx[127:96])
  );
AES_Comp_InvSubBytesComp  SB0 (
    .x({ dx[31:24], dx[55:48], dx[79:72], dx[103:96] }),
    .y(sb[31:0])
  );
AES_Comp_InvSubBytesComp  SB1 (
    .x({ dx[63:56], dx[87:80], dx[111:104], dx[7:0] }),
    .y(sb[63:32])
  );
AES_Comp_InvSubBytesComp  SB2 (
    .x({ dx[95:88], dx[119:112], dx[15:8], dx[39:32] }),
    .y(sb[95:64])
  );
AES_Comp_InvSubBytesComp  SB3 (
    .x({ dx[127:120], dx[23:16], dx[47:40], dx[71:64] }),
    .y(sb[127:96])
  );
AES_Comp_SubBytesComp  SBK (
    .x({ _068_, _067_, _065_, _064_, _063_, _062_, _061_, _060_, _059_, _058_, _057_, _056_, _054_, _053_, _052_, _051_, _050_, _049_, _048_, _047_, _046_, _045_, _075_, _074_, _073_, _072_, _071_, _070_, _069_, _066_, _055_, _044_ }),
    .y(so)
  );
assign  { _077_[5:2], _077_[0] } = { ki[60], ki[92], so[28], ki[124], Kgen };
assign  _081_[4:0] = { so[25], ki[121], ki[89], _078_[1], Kgen };
assign  { _076_[5:2], _076_[0] } = { ki[62], ki[94], so[30], ki[126], Kgen };
assign  { _015_[5:3], _015_[0] } = { so[27], ki[123], ki[91], Kgen };
assign  _079_[4:0] = { so[30], ki[126], ki[94], _076_[1], Kgen };
assign  _000_[6:1] = { so[24], ki[120], ki[88], Rrg[0], Kgen, Rrg[8] };
assign  { _078_[5:2], _078_[0] } = { ki[57], ki[89], so[25], ki[121], Kgen };
assign  { _025_[5:3], _025_[1:0] } = { so[31], ki[127], ki[95], _021_[2], Kgen };
assign  { _021_[5:3], _021_[0] } = { so[29], ki[125], ki[93], Kgen };
assign  { _011_[5:3], _011_[0] } = { so[26], ki[122], ki[90], Kgen };
assign  _080_[4:0] = { so[28], ki[124], ki[92], _077_[1], Kgen };
assign  \rcon$func$AES_Comp.v:408$441.x  = 10'hxxx;
assign  \rcon$func$AES_Comp.v:412$442.x  = 10'hxxx;
assign  sr = { dx[127:120], dx[23:16], dx[47:40], dx[71:64], dx[95:88], dx[119:112], dx[15:8], dx[39:32], dx[63:56], dx[87:80], dx[111:104], dx[7:0], dx[31:24], dx[55:48], dx[79:72], dx[103:96] };
endmodule
