module Trojan_Trigger(rst,  state, Tj_Trig);
wire  _000_;
wire  _001_;
wire  _002_;
wire  _003_;
wire  _004_;
wire  _005_;
wire  _006_;
wire  _007_;
wire  _008_;
wire  _009_;
wire  _010_;
wire  _011_;
wire  _012_;
wire  [7:0] _013_;
wire  _014_;
wire  _015_;
wire  _016_;
wire  _017_;
wire  _018_;
wire  _019_;
wire  _020_;
wire  _021_;
wire  _022_;
wire  _023_;
wire  _024_;
wire  _025_;
wire  _026_;
wire  _027_;
wire  _028_;
wire  _029_;
wire  _030_;
wire  _031_;
wire  _032_;
wire  _033_;
wire  _034_;
wire  _035_;
wire  _036_;
wire  _037_;
wire  _038_;
wire  _039_;
wire  _040_;
wire  _041_;
wire  [5:0] _042_;
wire  [5:0] _043_;
wire  [5:0] _044_;
wire  [5:0] _045_;
wire  [5:0] _046_;
output  Tj_Trig;
input  rst;
input  [127:0] state;
LUT6  #(
    .INIT(64'h000000007fffffff)
  ) _047_ (
    .I0(_046_[0]),
    .I1(_046_[1]),
    .I2(_046_[2]),
    .I3(_046_[3]),
    .I4(_046_[4]),
    .I5(rst),
    .O(_041_)
  );
LUT6  #(
    .INIT(64'h0001000000000000)
  ) _048_ (
    .I0(state[58]),
    .I1(state[60]),
    .I2(state[61]),
    .I3(state[62]),
    .I4(_042_[4]),
    .I5(_042_[5]),
    .O(_046_[4])
  );
LUT4  #(
    .INIT(16'h0001)
  ) _049_ (
    .I0(state[53]),
    .I1(state[54]),
    .I2(state[56]),
    .I3(state[57]),
    .O(_042_[4])
  );
LUT6  #(
    .INIT(64'h0000000000000001)
  ) _050_ (
    .I0(state[67]),
    .I1(state[71]),
    .I2(state[72]),
    .I3(state[75]),
    .I4(state[76]),
    .I5(state[79]),
    .O(_003_)
  );
MUXF7  _051_ (
    .I0(_003_),
    .I1(1'h0),
    .O(_001_),
    .S(state[81])
  );
MUXF7  _052_ (
    .I0(1'h0),
    .I1(1'h0),
    .O(_002_),
    .S(state[81])
  );
MUXF8  _053_ (
    .I0(_001_),
    .I1(_002_),
    .O(_042_[5]),
    .S(state[83])
  );
LUT6  #(
    .INIT(64'h0001000000000000)
  ) _054_ (
    .I0(state[24]),
    .I1(state[25]),
    .I2(state[28]),
    .I3(state[29]),
    .I4(_043_[4]),
    .I5(_043_[5]),
    .O(_046_[0])
  );
LUT4  #(
    .INIT(16'h0001)
  ) _055_ (
    .I0(state[8]),
    .I1(state[12]),
    .I2(state[17]),
    .I3(state[21]),
    .O(_043_[4])
  );
LUT6  #(
    .INIT(64'h0000000000000001)
  ) _056_ (
    .I0(state[34]),
    .I1(state[38]),
    .I2(state[40]),
    .I3(state[42]),
    .I4(state[44]),
    .I5(state[46]),
    .O(_006_)
  );
MUXF7  _057_ (
    .I0(_006_),
    .I1(1'h0),
    .O(_004_),
    .S(state[49])
  );
MUXF7  _058_ (
    .I0(1'h0),
    .I1(1'h0),
    .O(_005_),
    .S(state[49])
  );
MUXF8  _059_ (
    .I0(_004_),
    .I1(_005_),
    .O(_043_[5]),
    .S(state[50])
  );
LUT6  #(
    .INIT(64'h0001000000000000)
  ) _060_ (
    .I0(state[115]),
    .I1(state[117]),
    .I2(state[118]),
    .I3(state[119]),
    .I4(_044_[4]),
    .I5(_044_[5]),
    .O(_046_[1])
  );
LUT4  #(
    .INIT(16'h0001)
  ) _061_ (
    .I0(state[110]),
    .I1(state[111]),
    .I2(state[113]),
    .I3(state[114]),
    .O(_044_[4])
  );
LUT6  #(
    .INIT(64'h0000000000000001)
  ) _062_ (
    .I0(state[120]),
    .I1(state[121]),
    .I2(state[122]),
    .I3(state[123]),
    .I4(state[124]),
    .I5(state[125]),
    .O(_009_)
  );
MUXF7  _063_ (
    .I0(_009_),
    .I1(1'h0),
    .O(_007_),
    .S(state[126])
  );
MUXF7  _064_ (
    .I0(1'h0),
    .I1(1'h0),
    .O(_008_),
    .S(state[126])
  );
MUXF8  _065_ (
    .I0(_007_),
    .I1(_008_),
    .O(_044_[5]),
    .S(state[127])
  );
LUT6  #(
    .INIT(64'h0001000000000000)
  ) _066_ (
    .I0(state[91]),
    .I1(state[92]),
    .I2(state[93]),
    .I3(state[95]),
    .I4(_045_[4]),
    .I5(_045_[5]),
    .O(_046_[2])
  );
LUT4  #(
    .INIT(16'h0001)
  ) _067_ (
    .I0(state[85]),
    .I1(state[87]),
    .I2(state[88]),
    .I3(state[89]),
    .O(_045_[4])
  );
LUT6  #(
    .INIT(64'h0000000000000001)
  ) _068_ (
    .I0(state[98]),
    .I1(state[99]),
    .I2(state[102]),
    .I3(state[103]),
    .I4(state[104]),
    .I5(state[106]),
    .O(_012_)
  );
MUXF7  _069_ (
    .I0(_012_),
    .I1(1'h0),
    .O(_010_),
    .S(state[107])
  );
MUXF7  _070_ (
    .I0(1'h0),
    .I1(1'h0),
    .O(_011_),
    .S(state[107])
  );
MUXF8  _071_ (
    .I0(_010_),
    .I1(_011_),
    .O(_045_[5]),
    .S(state[108])
  );
MUXF7  _072_ (
    .I0(1'h0),
    .I1(1'h0),
    .O(_014_),
    .S(_013_[6])
  );
LUT6  #(
    .INIT(64'h8000000000000000)
  ) _073_ (
    .I0(_013_[0]),
    .I1(_013_[1]),
    .I2(_013_[2]),
    .I3(_013_[3]),
    .I4(_013_[4]),
    .I5(_013_[5]),
    .O(_016_)
  );
MUXF7  _074_ (
    .I0(1'h0),
    .I1(_016_),
    .O(_015_),
    .S(_013_[6])
  );
MUXF8  _075_ (
    .I0(_014_),
    .I1(_015_),
    .O(_046_[3]),
    .S(_013_[7])
  );
MUXF7  _076_ (
    .I0(1'h0),
    .I1(1'h0),
    .O(_017_),
    .S(state[30])
  );
LUT6  #(
    .INIT(64'h8000000000000000)
  ) _077_ (
    .I0(state[19]),
    .I1(state[20]),
    .I2(state[22]),
    .I3(state[23]),
    .I4(state[26]),
    .I5(state[27]),
    .O(_019_)
  );
MUXF7  _078_ (
    .I0(1'h0),
    .I1(_019_),
    .O(_018_),
    .S(state[30])
  );
MUXF8  _079_ (
    .I0(_017_),
    .I1(_018_),
    .O(_013_[0]),
    .S(state[31])
  );
MUXF7  _080_ (
    .I0(1'h0),
    .I1(1'h0),
    .O(_020_),
    .S(state[41])
  );
LUT6  #(
    .INIT(64'h8000000000000000)
  ) _081_ (
    .I0(state[32]),
    .I1(state[33]),
    .I2(state[35]),
    .I3(state[36]),
    .I4(state[37]),
    .I5(state[39]),
    .O(_022_)
  );
MUXF7  _082_ (
    .I0(1'h0),
    .I1(_022_),
    .O(_021_),
    .S(state[41])
  );
MUXF8  _083_ (
    .I0(_020_),
    .I1(_021_),
    .O(_013_[1]),
    .S(state[43])
  );
MUXF7  _084_ (
    .I0(1'h0),
    .I1(1'h0),
    .O(_023_),
    .S(state[6])
  );
LUT6  #(
    .INIT(64'h8000000000000000)
  ) _085_ (
    .I0(state[0]),
    .I1(state[1]),
    .I2(state[2]),
    .I3(state[3]),
    .I4(state[4]),
    .I5(state[5]),
    .O(_025_)
  );
MUXF7  _086_ (
    .I0(1'h0),
    .I1(_025_),
    .O(_024_),
    .S(state[6])
  );
MUXF8  _087_ (
    .I0(_023_),
    .I1(_024_),
    .O(_013_[2]),
    .S(state[7])
  );
MUXF7  _088_ (
    .I0(1'h0),
    .I1(1'h0),
    .O(_026_),
    .S(state[16])
  );
LUT6  #(
    .INIT(64'h8000000000000000)
  ) _089_ (
    .I0(state[9]),
    .I1(state[10]),
    .I2(state[11]),
    .I3(state[13]),
    .I4(state[14]),
    .I5(state[15]),
    .O(_028_)
  );
MUXF7  _090_ (
    .I0(1'h0),
    .I1(_028_),
    .O(_027_),
    .S(state[16])
  );
MUXF8  _091_ (
    .I0(_026_),
    .I1(_027_),
    .O(_013_[3]),
    .S(state[18])
  );
MUXF7  _092_ (
    .I0(1'h0),
    .I1(1'h0),
    .O(_029_),
    .S(state[90])
  );
LUT6  #(
    .INIT(64'h8000000000000000)
  ) _093_ (
    .I0(state[77]),
    .I1(state[78]),
    .I2(state[80]),
    .I3(state[82]),
    .I4(state[84]),
    .I5(state[86]),
    .O(_031_)
  );
MUXF7  _094_ (
    .I0(1'h0),
    .I1(_031_),
    .O(_030_),
    .S(state[90])
  );
MUXF8  _095_ (
    .I0(_029_),
    .I1(_030_),
    .O(_013_[4]),
    .S(state[94])
  );
MUXF7  _096_ (
    .I0(1'h0),
    .I1(1'h0),
    .O(_032_),
    .S(state[112])
  );
LUT6  #(
    .INIT(64'h8000000000000000)
  ) _097_ (
    .I0(state[96]),
    .I1(state[97]),
    .I2(state[100]),
    .I3(state[101]),
    .I4(state[105]),
    .I5(state[109]),
    .O(_034_)
  );
MUXF7  _098_ (
    .I0(1'h0),
    .I1(_034_),
    .O(_033_),
    .S(state[112])
  );
MUXF8  _099_ (
    .I0(_032_),
    .I1(_033_),
    .O(_013_[5]),
    .S(state[116])
  );
MUXF7  _100_ (
    .I0(1'h0),
    .I1(1'h0),
    .O(_035_),
    .S(state[59])
  );
LUT6  #(
    .INIT(64'h8000000000000000)
  ) _101_ (
    .I0(state[45]),
    .I1(state[47]),
    .I2(state[48]),
    .I3(state[51]),
    .I4(state[52]),
    .I5(state[55]),
    .O(_037_)
  );
MUXF7  _102_ (
    .I0(1'h0),
    .I1(_037_),
    .O(_036_),
    .S(state[59])
  );
MUXF8  _103_ (
    .I0(_035_),
    .I1(_036_),
    .O(_013_[6]),
    .S(state[63])
  );
MUXF7  _104_ (
    .I0(1'h0),
    .I1(1'h0),
    .O(_038_),
    .S(state[73])
  );
LUT6  #(
    .INIT(64'h8000000000000000)
  ) _105_ (
    .I0(state[64]),
    .I1(state[65]),
    .I2(state[66]),
    .I3(state[68]),
    .I4(state[69]),
    .I5(state[70]),
    .O(_040_)
  );
MUXF7  _106_ (
    .I0(1'h0),
    .I1(_040_),
    .O(_039_),
    .S(state[73])
  );
MUXF8  _107_ (
    .I0(_038_),
    .I1(_039_),
    .O(_013_[7]),
    .S(state[74])
  );
INV  _108_ (
    .I(rst),
    .O(_000_)
  );
LDCE  #(
    .INIT(1'hx),
    .IS_G_INVERTED(1'h1)
  ) _109_ (
    .CLR(1'h0),
    .D(_000_),
    .G(_041_),
    .GE(1'h1),
    .Q(Tj_Trig)
  );
assign  _043_[3:0] = { state[29:28], state[25:24] };
assign  _042_[3:0] = { state[62:60], state[58] };
assign  _046_[5] = rst;
assign  _045_[3:0] = { state[95], state[93:91] };
assign  _044_[3:0] = { state[119:117], state[115] };
endmodule
