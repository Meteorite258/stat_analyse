module final_round(clk,  state_in, key_in, state_out);
input  clk;
wire  [31:0] k0;
wire  [31:0] k1;
wire  [31:0] k2;
wire  [31:0] k3;
input  [127:0] key_in;
wire  [7:0] p00;
wire  [7:0] p01;
wire  [7:0] p02;
wire  [7:0] p03;
wire  [7:0] p10;
wire  [7:0] p11;
wire  [7:0] p12;
wire  [7:0] p13;
wire  [7:0] p20;
wire  [7:0] p21;
wire  [7:0] p22;
wire  [7:0] p23;
wire  [7:0] p30;
wire  [7:0] p31;
wire  [7:0] p32;
wire  [7:0] p33;
wire  [31:0] s0;
wire  [31:0] s1;
wire  [31:0] s2;
wire  [31:0] s3;
input  [127:0] state_in;
output  [127:0] state_out;
wire  [31:0] z0;
wire  [31:0] z1;
wire  [31:0] z2;
wire  [31:0] z3;
LUT2  #(
    .INIT(4'h6)
  ) _000_ (
    .I0(p33[0]),
    .I1(key_in[96]),
    .O(z0[0])
  );
LUT2  #(
    .INIT(4'h6)
  ) _001_ (
    .I0(p33[1]),
    .I1(key_in[97]),
    .O(z0[1])
  );
LUT2  #(
    .INIT(4'h6)
  ) _002_ (
    .I0(p33[2]),
    .I1(key_in[98]),
    .O(z0[2])
  );
LUT2  #(
    .INIT(4'h6)
  ) _003_ (
    .I0(p33[3]),
    .I1(key_in[99]),
    .O(z0[3])
  );
LUT2  #(
    .INIT(4'h6)
  ) _004_ (
    .I0(p33[4]),
    .I1(key_in[100]),
    .O(z0[4])
  );
LUT2  #(
    .INIT(4'h6)
  ) _005_ (
    .I0(p33[5]),
    .I1(key_in[101]),
    .O(z0[5])
  );
LUT2  #(
    .INIT(4'h6)
  ) _006_ (
    .I0(p33[6]),
    .I1(key_in[102]),
    .O(z0[6])
  );
LUT2  #(
    .INIT(4'h6)
  ) _007_ (
    .I0(p33[7]),
    .I1(key_in[103]),
    .O(z0[7])
  );
LUT2  #(
    .INIT(4'h6)
  ) _008_ (
    .I0(p22[0]),
    .I1(key_in[104]),
    .O(z0[8])
  );
LUT2  #(
    .INIT(4'h6)
  ) _009_ (
    .I0(p22[1]),
    .I1(key_in[105]),
    .O(z0[9])
  );
LUT2  #(
    .INIT(4'h6)
  ) _010_ (
    .I0(p22[2]),
    .I1(key_in[106]),
    .O(z0[10])
  );
LUT2  #(
    .INIT(4'h6)
  ) _011_ (
    .I0(p22[3]),
    .I1(key_in[107]),
    .O(z0[11])
  );
LUT2  #(
    .INIT(4'h6)
  ) _012_ (
    .I0(p22[4]),
    .I1(key_in[108]),
    .O(z0[12])
  );
LUT2  #(
    .INIT(4'h6)
  ) _013_ (
    .I0(p22[5]),
    .I1(key_in[109]),
    .O(z0[13])
  );
LUT2  #(
    .INIT(4'h6)
  ) _014_ (
    .I0(p22[6]),
    .I1(key_in[110]),
    .O(z0[14])
  );
LUT2  #(
    .INIT(4'h6)
  ) _015_ (
    .I0(p22[7]),
    .I1(key_in[111]),
    .O(z0[15])
  );
LUT2  #(
    .INIT(4'h6)
  ) _016_ (
    .I0(p11[0]),
    .I1(key_in[112]),
    .O(z0[16])
  );
LUT2  #(
    .INIT(4'h6)
  ) _017_ (
    .I0(p11[1]),
    .I1(key_in[113]),
    .O(z0[17])
  );
LUT2  #(
    .INIT(4'h6)
  ) _018_ (
    .I0(p11[2]),
    .I1(key_in[114]),
    .O(z0[18])
  );
LUT2  #(
    .INIT(4'h6)
  ) _019_ (
    .I0(p11[3]),
    .I1(key_in[115]),
    .O(z0[19])
  );
LUT2  #(
    .INIT(4'h6)
  ) _020_ (
    .I0(p11[4]),
    .I1(key_in[116]),
    .O(z0[20])
  );
LUT2  #(
    .INIT(4'h6)
  ) _021_ (
    .I0(p11[5]),
    .I1(key_in[117]),
    .O(z0[21])
  );
LUT2  #(
    .INIT(4'h6)
  ) _022_ (
    .I0(p11[6]),
    .I1(key_in[118]),
    .O(z0[22])
  );
LUT2  #(
    .INIT(4'h6)
  ) _023_ (
    .I0(p11[7]),
    .I1(key_in[119]),
    .O(z0[23])
  );
LUT2  #(
    .INIT(4'h6)
  ) _024_ (
    .I0(p00[0]),
    .I1(key_in[120]),
    .O(z0[24])
  );
LUT2  #(
    .INIT(4'h6)
  ) _025_ (
    .I0(p00[1]),
    .I1(key_in[121]),
    .O(z0[25])
  );
LUT2  #(
    .INIT(4'h6)
  ) _026_ (
    .I0(p00[2]),
    .I1(key_in[122]),
    .O(z0[26])
  );
LUT2  #(
    .INIT(4'h6)
  ) _027_ (
    .I0(p00[3]),
    .I1(key_in[123]),
    .O(z0[27])
  );
LUT2  #(
    .INIT(4'h6)
  ) _028_ (
    .I0(p00[4]),
    .I1(key_in[124]),
    .O(z0[28])
  );
LUT2  #(
    .INIT(4'h6)
  ) _029_ (
    .I0(p00[5]),
    .I1(key_in[125]),
    .O(z0[29])
  );
LUT2  #(
    .INIT(4'h6)
  ) _030_ (
    .I0(p00[6]),
    .I1(key_in[126]),
    .O(z0[30])
  );
LUT2  #(
    .INIT(4'h6)
  ) _031_ (
    .I0(p00[7]),
    .I1(key_in[127]),
    .O(z0[31])
  );
LUT2  #(
    .INIT(4'h6)
  ) _032_ (
    .I0(p03[0]),
    .I1(key_in[64]),
    .O(z1[0])
  );
LUT2  #(
    .INIT(4'h6)
  ) _033_ (
    .I0(p03[1]),
    .I1(key_in[65]),
    .O(z1[1])
  );
LUT2  #(
    .INIT(4'h6)
  ) _034_ (
    .I0(p03[2]),
    .I1(key_in[66]),
    .O(z1[2])
  );
LUT2  #(
    .INIT(4'h6)
  ) _035_ (
    .I0(p03[3]),
    .I1(key_in[67]),
    .O(z1[3])
  );
LUT2  #(
    .INIT(4'h6)
  ) _036_ (
    .I0(p03[4]),
    .I1(key_in[68]),
    .O(z1[4])
  );
LUT2  #(
    .INIT(4'h6)
  ) _037_ (
    .I0(p03[5]),
    .I1(key_in[69]),
    .O(z1[5])
  );
LUT2  #(
    .INIT(4'h6)
  ) _038_ (
    .I0(p03[6]),
    .I1(key_in[70]),
    .O(z1[6])
  );
LUT2  #(
    .INIT(4'h6)
  ) _039_ (
    .I0(p03[7]),
    .I1(key_in[71]),
    .O(z1[7])
  );
LUT2  #(
    .INIT(4'h6)
  ) _040_ (
    .I0(p32[0]),
    .I1(key_in[72]),
    .O(z1[8])
  );
LUT2  #(
    .INIT(4'h6)
  ) _041_ (
    .I0(p32[1]),
    .I1(key_in[73]),
    .O(z1[9])
  );
LUT2  #(
    .INIT(4'h6)
  ) _042_ (
    .I0(p32[2]),
    .I1(key_in[74]),
    .O(z1[10])
  );
LUT2  #(
    .INIT(4'h6)
  ) _043_ (
    .I0(p32[3]),
    .I1(key_in[75]),
    .O(z1[11])
  );
LUT2  #(
    .INIT(4'h6)
  ) _044_ (
    .I0(p32[4]),
    .I1(key_in[76]),
    .O(z1[12])
  );
LUT2  #(
    .INIT(4'h6)
  ) _045_ (
    .I0(p32[5]),
    .I1(key_in[77]),
    .O(z1[13])
  );
LUT2  #(
    .INIT(4'h6)
  ) _046_ (
    .I0(p32[6]),
    .I1(key_in[78]),
    .O(z1[14])
  );
LUT2  #(
    .INIT(4'h6)
  ) _047_ (
    .I0(p32[7]),
    .I1(key_in[79]),
    .O(z1[15])
  );
LUT2  #(
    .INIT(4'h6)
  ) _048_ (
    .I0(p21[0]),
    .I1(key_in[80]),
    .O(z1[16])
  );
LUT2  #(
    .INIT(4'h6)
  ) _049_ (
    .I0(p21[1]),
    .I1(key_in[81]),
    .O(z1[17])
  );
LUT2  #(
    .INIT(4'h6)
  ) _050_ (
    .I0(p21[2]),
    .I1(key_in[82]),
    .O(z1[18])
  );
LUT2  #(
    .INIT(4'h6)
  ) _051_ (
    .I0(p21[3]),
    .I1(key_in[83]),
    .O(z1[19])
  );
LUT2  #(
    .INIT(4'h6)
  ) _052_ (
    .I0(p21[4]),
    .I1(key_in[84]),
    .O(z1[20])
  );
LUT2  #(
    .INIT(4'h6)
  ) _053_ (
    .I0(p21[5]),
    .I1(key_in[85]),
    .O(z1[21])
  );
LUT2  #(
    .INIT(4'h6)
  ) _054_ (
    .I0(p21[6]),
    .I1(key_in[86]),
    .O(z1[22])
  );
LUT2  #(
    .INIT(4'h6)
  ) _055_ (
    .I0(p21[7]),
    .I1(key_in[87]),
    .O(z1[23])
  );
LUT2  #(
    .INIT(4'h6)
  ) _056_ (
    .I0(p10[0]),
    .I1(key_in[88]),
    .O(z1[24])
  );
LUT2  #(
    .INIT(4'h6)
  ) _057_ (
    .I0(p10[1]),
    .I1(key_in[89]),
    .O(z1[25])
  );
LUT2  #(
    .INIT(4'h6)
  ) _058_ (
    .I0(p10[2]),
    .I1(key_in[90]),
    .O(z1[26])
  );
LUT2  #(
    .INIT(4'h6)
  ) _059_ (
    .I0(p10[3]),
    .I1(key_in[91]),
    .O(z1[27])
  );
LUT2  #(
    .INIT(4'h6)
  ) _060_ (
    .I0(p10[4]),
    .I1(key_in[92]),
    .O(z1[28])
  );
LUT2  #(
    .INIT(4'h6)
  ) _061_ (
    .I0(p10[5]),
    .I1(key_in[93]),
    .O(z1[29])
  );
LUT2  #(
    .INIT(4'h6)
  ) _062_ (
    .I0(p10[6]),
    .I1(key_in[94]),
    .O(z1[30])
  );
LUT2  #(
    .INIT(4'h6)
  ) _063_ (
    .I0(p10[7]),
    .I1(key_in[95]),
    .O(z1[31])
  );
LUT2  #(
    .INIT(4'h6)
  ) _064_ (
    .I0(p13[0]),
    .I1(key_in[32]),
    .O(z2[0])
  );
LUT2  #(
    .INIT(4'h6)
  ) _065_ (
    .I0(p13[1]),
    .I1(key_in[33]),
    .O(z2[1])
  );
LUT2  #(
    .INIT(4'h6)
  ) _066_ (
    .I0(p13[2]),
    .I1(key_in[34]),
    .O(z2[2])
  );
LUT2  #(
    .INIT(4'h6)
  ) _067_ (
    .I0(p13[3]),
    .I1(key_in[35]),
    .O(z2[3])
  );
LUT2  #(
    .INIT(4'h6)
  ) _068_ (
    .I0(p13[4]),
    .I1(key_in[36]),
    .O(z2[4])
  );
LUT2  #(
    .INIT(4'h6)
  ) _069_ (
    .I0(p13[5]),
    .I1(key_in[37]),
    .O(z2[5])
  );
LUT2  #(
    .INIT(4'h6)
  ) _070_ (
    .I0(p13[6]),
    .I1(key_in[38]),
    .O(z2[6])
  );
LUT2  #(
    .INIT(4'h6)
  ) _071_ (
    .I0(p13[7]),
    .I1(key_in[39]),
    .O(z2[7])
  );
LUT2  #(
    .INIT(4'h6)
  ) _072_ (
    .I0(p02[0]),
    .I1(key_in[40]),
    .O(z2[8])
  );
LUT2  #(
    .INIT(4'h6)
  ) _073_ (
    .I0(p02[1]),
    .I1(key_in[41]),
    .O(z2[9])
  );
LUT2  #(
    .INIT(4'h6)
  ) _074_ (
    .I0(p02[2]),
    .I1(key_in[42]),
    .O(z2[10])
  );
LUT2  #(
    .INIT(4'h6)
  ) _075_ (
    .I0(p02[3]),
    .I1(key_in[43]),
    .O(z2[11])
  );
LUT2  #(
    .INIT(4'h6)
  ) _076_ (
    .I0(p02[4]),
    .I1(key_in[44]),
    .O(z2[12])
  );
LUT2  #(
    .INIT(4'h6)
  ) _077_ (
    .I0(p02[5]),
    .I1(key_in[45]),
    .O(z2[13])
  );
LUT2  #(
    .INIT(4'h6)
  ) _078_ (
    .I0(p02[6]),
    .I1(key_in[46]),
    .O(z2[14])
  );
LUT2  #(
    .INIT(4'h6)
  ) _079_ (
    .I0(p02[7]),
    .I1(key_in[47]),
    .O(z2[15])
  );
LUT2  #(
    .INIT(4'h6)
  ) _080_ (
    .I0(p31[0]),
    .I1(key_in[48]),
    .O(z2[16])
  );
LUT2  #(
    .INIT(4'h6)
  ) _081_ (
    .I0(p31[1]),
    .I1(key_in[49]),
    .O(z2[17])
  );
LUT2  #(
    .INIT(4'h6)
  ) _082_ (
    .I0(p31[2]),
    .I1(key_in[50]),
    .O(z2[18])
  );
LUT2  #(
    .INIT(4'h6)
  ) _083_ (
    .I0(p31[3]),
    .I1(key_in[51]),
    .O(z2[19])
  );
LUT2  #(
    .INIT(4'h6)
  ) _084_ (
    .I0(p31[4]),
    .I1(key_in[52]),
    .O(z2[20])
  );
LUT2  #(
    .INIT(4'h6)
  ) _085_ (
    .I0(p31[5]),
    .I1(key_in[53]),
    .O(z2[21])
  );
LUT2  #(
    .INIT(4'h6)
  ) _086_ (
    .I0(p31[6]),
    .I1(key_in[54]),
    .O(z2[22])
  );
LUT2  #(
    .INIT(4'h6)
  ) _087_ (
    .I0(p31[7]),
    .I1(key_in[55]),
    .O(z2[23])
  );
LUT2  #(
    .INIT(4'h6)
  ) _088_ (
    .I0(p20[0]),
    .I1(key_in[56]),
    .O(z2[24])
  );
LUT2  #(
    .INIT(4'h6)
  ) _089_ (
    .I0(p20[1]),
    .I1(key_in[57]),
    .O(z2[25])
  );
LUT2  #(
    .INIT(4'h6)
  ) _090_ (
    .I0(p20[2]),
    .I1(key_in[58]),
    .O(z2[26])
  );
LUT2  #(
    .INIT(4'h6)
  ) _091_ (
    .I0(p20[3]),
    .I1(key_in[59]),
    .O(z2[27])
  );
LUT2  #(
    .INIT(4'h6)
  ) _092_ (
    .I0(p20[4]),
    .I1(key_in[60]),
    .O(z2[28])
  );
LUT2  #(
    .INIT(4'h6)
  ) _093_ (
    .I0(p20[5]),
    .I1(key_in[61]),
    .O(z2[29])
  );
LUT2  #(
    .INIT(4'h6)
  ) _094_ (
    .I0(p20[6]),
    .I1(key_in[62]),
    .O(z2[30])
  );
LUT2  #(
    .INIT(4'h6)
  ) _095_ (
    .I0(p20[7]),
    .I1(key_in[63]),
    .O(z2[31])
  );
LUT2  #(
    .INIT(4'h6)
  ) _096_ (
    .I0(p23[0]),
    .I1(key_in[0]),
    .O(z3[0])
  );
LUT2  #(
    .INIT(4'h6)
  ) _097_ (
    .I0(p23[1]),
    .I1(key_in[1]),
    .O(z3[1])
  );
LUT2  #(
    .INIT(4'h6)
  ) _098_ (
    .I0(p23[2]),
    .I1(key_in[2]),
    .O(z3[2])
  );
LUT2  #(
    .INIT(4'h6)
  ) _099_ (
    .I0(p23[3]),
    .I1(key_in[3]),
    .O(z3[3])
  );
LUT2  #(
    .INIT(4'h6)
  ) _100_ (
    .I0(p23[4]),
    .I1(key_in[4]),
    .O(z3[4])
  );
LUT2  #(
    .INIT(4'h6)
  ) _101_ (
    .I0(p23[5]),
    .I1(key_in[5]),
    .O(z3[5])
  );
LUT2  #(
    .INIT(4'h6)
  ) _102_ (
    .I0(p23[6]),
    .I1(key_in[6]),
    .O(z3[6])
  );
LUT2  #(
    .INIT(4'h6)
  ) _103_ (
    .I0(p23[7]),
    .I1(key_in[7]),
    .O(z3[7])
  );
LUT2  #(
    .INIT(4'h6)
  ) _104_ (
    .I0(p12[0]),
    .I1(key_in[8]),
    .O(z3[8])
  );
LUT2  #(
    .INIT(4'h6)
  ) _105_ (
    .I0(p12[1]),
    .I1(key_in[9]),
    .O(z3[9])
  );
LUT2  #(
    .INIT(4'h6)
  ) _106_ (
    .I0(p12[2]),
    .I1(key_in[10]),
    .O(z3[10])
  );
LUT2  #(
    .INIT(4'h6)
  ) _107_ (
    .I0(p12[3]),
    .I1(key_in[11]),
    .O(z3[11])
  );
LUT2  #(
    .INIT(4'h6)
  ) _108_ (
    .I0(p12[4]),
    .I1(key_in[12]),
    .O(z3[12])
  );
LUT2  #(
    .INIT(4'h6)
  ) _109_ (
    .I0(p12[5]),
    .I1(key_in[13]),
    .O(z3[13])
  );
LUT2  #(
    .INIT(4'h6)
  ) _110_ (
    .I0(p12[6]),
    .I1(key_in[14]),
    .O(z3[14])
  );
LUT2  #(
    .INIT(4'h6)
  ) _111_ (
    .I0(p12[7]),
    .I1(key_in[15]),
    .O(z3[15])
  );
LUT2  #(
    .INIT(4'h6)
  ) _112_ (
    .I0(p01[0]),
    .I1(key_in[16]),
    .O(z3[16])
  );
LUT2  #(
    .INIT(4'h6)
  ) _113_ (
    .I0(p01[1]),
    .I1(key_in[17]),
    .O(z3[17])
  );
LUT2  #(
    .INIT(4'h6)
  ) _114_ (
    .I0(p01[2]),
    .I1(key_in[18]),
    .O(z3[18])
  );
LUT2  #(
    .INIT(4'h6)
  ) _115_ (
    .I0(p01[3]),
    .I1(key_in[19]),
    .O(z3[19])
  );
LUT2  #(
    .INIT(4'h6)
  ) _116_ (
    .I0(p01[4]),
    .I1(key_in[20]),
    .O(z3[20])
  );
LUT2  #(
    .INIT(4'h6)
  ) _117_ (
    .I0(p01[5]),
    .I1(key_in[21]),
    .O(z3[21])
  );
LUT2  #(
    .INIT(4'h6)
  ) _118_ (
    .I0(p01[6]),
    .I1(key_in[22]),
    .O(z3[22])
  );
LUT2  #(
    .INIT(4'h6)
  ) _119_ (
    .I0(p01[7]),
    .I1(key_in[23]),
    .O(z3[23])
  );
LUT2  #(
    .INIT(4'h6)
  ) _120_ (
    .I0(p30[0]),
    .I1(key_in[24]),
    .O(z3[24])
  );
LUT2  #(
    .INIT(4'h6)
  ) _121_ (
    .I0(p30[1]),
    .I1(key_in[25]),
    .O(z3[25])
  );
LUT2  #(
    .INIT(4'h6)
  ) _122_ (
    .I0(p30[2]),
    .I1(key_in[26]),
    .O(z3[26])
  );
LUT2  #(
    .INIT(4'h6)
  ) _123_ (
    .I0(p30[3]),
    .I1(key_in[27]),
    .O(z3[27])
  );
LUT2  #(
    .INIT(4'h6)
  ) _124_ (
    .I0(p30[4]),
    .I1(key_in[28]),
    .O(z3[28])
  );
LUT2  #(
    .INIT(4'h6)
  ) _125_ (
    .I0(p30[5]),
    .I1(key_in[29]),
    .O(z3[29])
  );
LUT2  #(
    .INIT(4'h6)
  ) _126_ (
    .I0(p30[6]),
    .I1(key_in[30]),
    .O(z3[30])
  );
LUT2  #(
    .INIT(4'h6)
  ) _127_ (
    .I0(p30[7]),
    .I1(key_in[31]),
    .O(z3[31])
  );
FDRE  #(
    .INIT(1'hx)
  ) _128_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[0]),
    .Q(state_out[0]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _129_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[1]),
    .Q(state_out[1]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _130_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[2]),
    .Q(state_out[2]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _131_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[3]),
    .Q(state_out[3]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _132_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[4]),
    .Q(state_out[4]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _133_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[5]),
    .Q(state_out[5]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _134_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[6]),
    .Q(state_out[6]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _135_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[7]),
    .Q(state_out[7]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _136_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[8]),
    .Q(state_out[8]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _137_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[9]),
    .Q(state_out[9]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _138_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[10]),
    .Q(state_out[10]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _139_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[11]),
    .Q(state_out[11]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _140_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[12]),
    .Q(state_out[12]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _141_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[13]),
    .Q(state_out[13]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _142_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[14]),
    .Q(state_out[14]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _143_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[15]),
    .Q(state_out[15]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _144_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[16]),
    .Q(state_out[16]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _145_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[17]),
    .Q(state_out[17]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _146_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[18]),
    .Q(state_out[18]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _147_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[19]),
    .Q(state_out[19]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _148_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[20]),
    .Q(state_out[20]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _149_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[21]),
    .Q(state_out[21]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _150_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[22]),
    .Q(state_out[22]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _151_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[23]),
    .Q(state_out[23]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _152_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[24]),
    .Q(state_out[24]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _153_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[25]),
    .Q(state_out[25]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _154_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[26]),
    .Q(state_out[26]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _155_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[27]),
    .Q(state_out[27]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _156_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[28]),
    .Q(state_out[28]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _157_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[29]),
    .Q(state_out[29]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _158_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[30]),
    .Q(state_out[30]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _159_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[31]),
    .Q(state_out[31]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _160_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[0]),
    .Q(state_out[32]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _161_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[1]),
    .Q(state_out[33]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _162_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[2]),
    .Q(state_out[34]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _163_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[3]),
    .Q(state_out[35]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _164_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[4]),
    .Q(state_out[36]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _165_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[5]),
    .Q(state_out[37]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _166_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[6]),
    .Q(state_out[38]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _167_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[7]),
    .Q(state_out[39]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _168_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[8]),
    .Q(state_out[40]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _169_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[9]),
    .Q(state_out[41]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _170_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[10]),
    .Q(state_out[42]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _171_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[11]),
    .Q(state_out[43]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _172_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[12]),
    .Q(state_out[44]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _173_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[13]),
    .Q(state_out[45]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _174_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[14]),
    .Q(state_out[46]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _175_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[15]),
    .Q(state_out[47]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _176_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[16]),
    .Q(state_out[48]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _177_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[17]),
    .Q(state_out[49]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _178_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[18]),
    .Q(state_out[50]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _179_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[19]),
    .Q(state_out[51]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _180_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[20]),
    .Q(state_out[52]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _181_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[21]),
    .Q(state_out[53]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _182_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[22]),
    .Q(state_out[54]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _183_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[23]),
    .Q(state_out[55]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _184_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[24]),
    .Q(state_out[56]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _185_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[25]),
    .Q(state_out[57]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _186_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[26]),
    .Q(state_out[58]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _187_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[27]),
    .Q(state_out[59]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _188_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[28]),
    .Q(state_out[60]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _189_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[29]),
    .Q(state_out[61]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _190_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[30]),
    .Q(state_out[62]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _191_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[31]),
    .Q(state_out[63]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _192_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[0]),
    .Q(state_out[64]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _193_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[1]),
    .Q(state_out[65]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _194_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[2]),
    .Q(state_out[66]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _195_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[3]),
    .Q(state_out[67]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _196_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[4]),
    .Q(state_out[68]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _197_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[5]),
    .Q(state_out[69]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _198_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[6]),
    .Q(state_out[70]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _199_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[7]),
    .Q(state_out[71]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _200_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[8]),
    .Q(state_out[72]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _201_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[9]),
    .Q(state_out[73]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _202_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[10]),
    .Q(state_out[74]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _203_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[11]),
    .Q(state_out[75]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _204_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[12]),
    .Q(state_out[76]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _205_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[13]),
    .Q(state_out[77]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _206_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[14]),
    .Q(state_out[78]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _207_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[15]),
    .Q(state_out[79]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _208_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[16]),
    .Q(state_out[80]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _209_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[17]),
    .Q(state_out[81]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _210_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[18]),
    .Q(state_out[82]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _211_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[19]),
    .Q(state_out[83]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _212_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[20]),
    .Q(state_out[84]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _213_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[21]),
    .Q(state_out[85]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _214_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[22]),
    .Q(state_out[86]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _215_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[23]),
    .Q(state_out[87]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _216_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[24]),
    .Q(state_out[88]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _217_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[25]),
    .Q(state_out[89]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _218_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[26]),
    .Q(state_out[90]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _219_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[27]),
    .Q(state_out[91]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _220_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[28]),
    .Q(state_out[92]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _221_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[29]),
    .Q(state_out[93]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _222_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[30]),
    .Q(state_out[94]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _223_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[31]),
    .Q(state_out[95]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _224_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[0]),
    .Q(state_out[96]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _225_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[1]),
    .Q(state_out[97]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _226_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[2]),
    .Q(state_out[98]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _227_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[3]),
    .Q(state_out[99]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _228_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[4]),
    .Q(state_out[100]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _229_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[5]),
    .Q(state_out[101]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _230_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[6]),
    .Q(state_out[102]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _231_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[7]),
    .Q(state_out[103]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _232_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[8]),
    .Q(state_out[104]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _233_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[9]),
    .Q(state_out[105]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _234_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[10]),
    .Q(state_out[106]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _235_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[11]),
    .Q(state_out[107]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _236_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[12]),
    .Q(state_out[108]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _237_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[13]),
    .Q(state_out[109]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _238_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[14]),
    .Q(state_out[110]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _239_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[15]),
    .Q(state_out[111]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _240_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[16]),
    .Q(state_out[112]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _241_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[17]),
    .Q(state_out[113]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _242_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[18]),
    .Q(state_out[114]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _243_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[19]),
    .Q(state_out[115]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _244_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[20]),
    .Q(state_out[116]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _245_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[21]),
    .Q(state_out[117]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _246_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[22]),
    .Q(state_out[118]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _247_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[23]),
    .Q(state_out[119]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _248_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[24]),
    .Q(state_out[120]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _249_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[25]),
    .Q(state_out[121]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _250_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[26]),
    .Q(state_out[122]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _251_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[27]),
    .Q(state_out[123]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _252_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[28]),
    .Q(state_out[124]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _253_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[29]),
    .Q(state_out[125]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _254_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[30]),
    .Q(state_out[126]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _255_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[31]),
    .Q(state_out[127]),
    .R(1'h0)
  );
S4  S4_1 (
    .clk(clk),
    .in(state_in[127:96]),
    .out({ p00, p01, p02, p03 })
  );
S4  S4_2 (
    .clk(clk),
    .in(state_in[95:64]),
    .out({ p10, p11, p12, p13 })
  );
S4  S4_3 (
    .clk(clk),
    .in(state_in[63:32]),
    .out({ p20, p21, p22, p23 })
  );
S4  S4_4 (
    .clk(clk),
    .in(state_in[31:0]),
    .out({ p30, p31, p32, p33 })
  );
assign  k0 = key_in[127:96];
assign  k1 = key_in[95:64];
assign  k2 = key_in[63:32];
assign  k3 = key_in[31:0];
assign  s0 = state_in[127:96];
assign  s1 = state_in[95:64];
assign  s2 = state_in[63:32];
assign  s3 = state_in[31:0];
endmodule
