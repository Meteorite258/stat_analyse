module AES_Comp(Kin,  Din, Dout, Krdy, Drdy, EncDec, RSTn, EN, CLK, BSY, Kvld, Dvld);
wire  _000_;
wire  _001_;
wire  _002_;
wire  _003_;
wire  _004_;
wire  _005_;
wire  _006_;
wire  _007_;
wire  _008_;
wire  _009_;
wire  _010_;
wire  _011_;
wire  _012_;
wire  _013_;
wire  _014_;
wire  _015_;
wire  _016_;
wire  _017_;
wire  _018_;
wire  _019_;
wire  _020_;
wire  _021_;
wire  _022_;
wire  _023_;
wire  _024_;
wire  _025_;
wire  _026_;
wire  _027_;
wire  _028_;
wire  _029_;
wire  _030_;
wire  _031_;
wire  _032_;
wire  _033_;
wire  _034_;
wire  _035_;
wire  _036_;
wire  _037_;
wire  _038_;
wire  _039_;
wire  _040_;
wire  _041_;
wire  _042_;
wire  _043_;
wire  _044_;
wire  _045_;
wire  _046_;
wire  _047_;
wire  _048_;
wire  _049_;
wire  _050_;
wire  _051_;
wire  _052_;
wire  _053_;
wire  _054_;
wire  _055_;
wire  _056_;
wire  _057_;
wire  _058_;
wire  _059_;
wire  _060_;
wire  _061_;
wire  _062_;
wire  _063_;
wire  _064_;
wire  _065_;
wire  _066_;
wire  _067_;
wire  _068_;
wire  _069_;
wire  _070_;
wire  _071_;
wire  _072_;
wire  _073_;
wire  _074_;
wire  _075_;
wire  _076_;
wire  _077_;
wire  _078_;
wire  _079_;
wire  _080_;
wire  _081_;
wire  _082_;
wire  _083_;
wire  _084_;
wire  _085_;
wire  _086_;
wire  _087_;
wire  _088_;
wire  _089_;
wire  _090_;
wire  _091_;
wire  _092_;
wire  _093_;
wire  _094_;
wire  _095_;
wire  _096_;
wire  _097_;
wire  _098_;
wire  _099_;
wire  _100_;
wire  _101_;
wire  _102_;
wire  _103_;
wire  _104_;
wire  _105_;
wire  _106_;
wire  _107_;
wire  _108_;
wire  _109_;
wire  _110_;
wire  _111_;
wire  _112_;
wire  _113_;
wire  _114_;
wire  _115_;
wire  _116_;
wire  _117_;
wire  _118_;
wire  _119_;
wire  _120_;
wire  _121_;
wire  _122_;
wire  _123_;
wire  _124_;
wire  _125_;
wire  _126_;
wire  _127_;
wire  _128_;
wire  _129_;
wire  _130_;
wire  _131_;
wire  _132_;
wire  _133_;
wire  _134_;
wire  [127:0] _135_;
wire  _136_;
wire  [127:0] _137_;
wire  _138_;
wire  _139_;
wire  [1:0] _140_;
output  BSY;
wire  BSY;
wire  BSY_D;
wire  BSY_E;
input  CLK;
wire  CLK;
input  [127:0] Din;
wire  [127:0] Din;
output  [127:0] Dout;
wire  [127:0] Dout;
wire  [127:0] Dout_D;
wire  [127:0] Dout_E;
input  Drdy;
wire  Drdy;
output  Dvld;
wire  Dvld;
wire  Dvld_D;
wire  Dvld_E;
wire  Dvld_reg;
input  EN;
wire  EN;
wire  EN_D;
wire  EN_E;
input  EncDec;
wire  EncDec;
input  [127:0] Kin;
wire  [127:0] Kin;
input  Krdy;
wire  Krdy;
output  Kvld;
wire  Kvld;
wire  Kvld_D;
wire  Kvld_E;
wire  Kvld_reg;
input  RSTn;
wire  RSTn;
LUT4  #(
    .INIT(16'h0c0a)
  ) _141_ (
    .I0(Dvld_E),
    .I1(Dvld_D),
    .I2(Dvld_reg),
    .I3(_140_[0]),
    .O(_129_)
  );
LUT4  #(
    .INIT(16'h0c0a)
  ) _142_ (
    .I0(Kvld_E),
    .I1(Kvld_D),
    .I2(Kvld_reg),
    .I3(_140_[0]),
    .O(_130_)
  );
LUT3  #(
    .INIT(8'hac)
  ) _143_ (
    .I0(Dout_D[0]),
    .I1(Dout_E[0]),
    .I2(_140_[0]),
    .O(_001_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _144_ (
    .I0(Dout_E[1]),
    .I1(Dout_D[1]),
    .I2(_140_[0]),
    .O(_040_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _145_ (
    .I0(Dout_E[2]),
    .I1(Dout_D[2]),
    .I2(_140_[0]),
    .O(_051_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _146_ (
    .I0(Dout_E[3]),
    .I1(Dout_D[3]),
    .I2(_140_[0]),
    .O(_062_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _147_ (
    .I0(Dout_E[4]),
    .I1(Dout_D[4]),
    .I2(_140_[0]),
    .O(_073_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _148_ (
    .I0(Dout_E[5]),
    .I1(Dout_D[5]),
    .I2(_140_[0]),
    .O(_084_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _149_ (
    .I0(Dout_E[6]),
    .I1(Dout_D[6]),
    .I2(_140_[0]),
    .O(_095_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _150_ (
    .I0(Dout_E[7]),
    .I1(Dout_D[7]),
    .I2(_140_[0]),
    .O(_106_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _151_ (
    .I0(Dout_E[8]),
    .I1(Dout_D[8]),
    .I2(_140_[0]),
    .O(_117_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _152_ (
    .I0(Dout_E[9]),
    .I1(Dout_D[9]),
    .I2(_140_[0]),
    .O(_128_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _153_ (
    .I0(Dout_E[10]),
    .I1(Dout_D[10]),
    .I2(_140_[0]),
    .O(_012_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _154_ (
    .I0(Dout_E[11]),
    .I1(Dout_D[11]),
    .I2(_140_[0]),
    .O(_023_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _155_ (
    .I0(Dout_E[12]),
    .I1(Dout_D[12]),
    .I2(_140_[0]),
    .O(_032_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _156_ (
    .I0(Dout_E[13]),
    .I1(Dout_D[13]),
    .I2(_140_[0]),
    .O(_033_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _157_ (
    .I0(Dout_E[14]),
    .I1(Dout_D[14]),
    .I2(_140_[0]),
    .O(_034_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _158_ (
    .I0(Dout_E[15]),
    .I1(Dout_D[15]),
    .I2(_140_[0]),
    .O(_035_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _159_ (
    .I0(Dout_E[16]),
    .I1(Dout_D[16]),
    .I2(_140_[0]),
    .O(_036_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _160_ (
    .I0(Dout_E[17]),
    .I1(Dout_D[17]),
    .I2(_140_[0]),
    .O(_037_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _161_ (
    .I0(Dout_E[18]),
    .I1(Dout_D[18]),
    .I2(_140_[0]),
    .O(_038_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _162_ (
    .I0(Dout_E[19]),
    .I1(Dout_D[19]),
    .I2(_140_[0]),
    .O(_039_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _163_ (
    .I0(Dout_E[20]),
    .I1(Dout_D[20]),
    .I2(_140_[0]),
    .O(_041_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _164_ (
    .I0(Dout_E[21]),
    .I1(Dout_D[21]),
    .I2(_140_[0]),
    .O(_042_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _165_ (
    .I0(Dout_E[22]),
    .I1(Dout_D[22]),
    .I2(_140_[0]),
    .O(_043_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _166_ (
    .I0(Dout_E[23]),
    .I1(Dout_D[23]),
    .I2(_140_[0]),
    .O(_044_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _167_ (
    .I0(Dout_E[24]),
    .I1(Dout_D[24]),
    .I2(_140_[0]),
    .O(_045_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _168_ (
    .I0(Dout_E[25]),
    .I1(Dout_D[25]),
    .I2(_140_[0]),
    .O(_046_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _169_ (
    .I0(Dout_E[26]),
    .I1(Dout_D[26]),
    .I2(_140_[0]),
    .O(_047_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _170_ (
    .I0(Dout_E[27]),
    .I1(Dout_D[27]),
    .I2(_140_[0]),
    .O(_048_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _171_ (
    .I0(Dout_E[28]),
    .I1(Dout_D[28]),
    .I2(_140_[0]),
    .O(_049_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _172_ (
    .I0(Dout_E[29]),
    .I1(Dout_D[29]),
    .I2(_140_[0]),
    .O(_050_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _173_ (
    .I0(Dout_E[30]),
    .I1(Dout_D[30]),
    .I2(_140_[0]),
    .O(_052_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _174_ (
    .I0(Dout_E[31]),
    .I1(Dout_D[31]),
    .I2(_140_[0]),
    .O(_053_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _175_ (
    .I0(Dout_E[32]),
    .I1(Dout_D[32]),
    .I2(_140_[0]),
    .O(_054_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _176_ (
    .I0(Dout_E[33]),
    .I1(Dout_D[33]),
    .I2(_140_[0]),
    .O(_055_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _177_ (
    .I0(Dout_E[34]),
    .I1(Dout_D[34]),
    .I2(_140_[0]),
    .O(_056_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _178_ (
    .I0(Dout_E[35]),
    .I1(Dout_D[35]),
    .I2(_140_[0]),
    .O(_057_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _179_ (
    .I0(Dout_E[36]),
    .I1(Dout_D[36]),
    .I2(_140_[0]),
    .O(_058_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _180_ (
    .I0(Dout_E[37]),
    .I1(Dout_D[37]),
    .I2(_140_[0]),
    .O(_059_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _181_ (
    .I0(Dout_E[38]),
    .I1(Dout_D[38]),
    .I2(_140_[0]),
    .O(_060_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _182_ (
    .I0(Dout_E[39]),
    .I1(Dout_D[39]),
    .I2(_140_[0]),
    .O(_061_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _183_ (
    .I0(Dout_E[40]),
    .I1(Dout_D[40]),
    .I2(_140_[0]),
    .O(_063_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _184_ (
    .I0(Dout_E[41]),
    .I1(Dout_D[41]),
    .I2(_140_[0]),
    .O(_064_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _185_ (
    .I0(Dout_E[42]),
    .I1(Dout_D[42]),
    .I2(_140_[0]),
    .O(_065_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _186_ (
    .I0(Dout_E[43]),
    .I1(Dout_D[43]),
    .I2(_140_[0]),
    .O(_066_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _187_ (
    .I0(Dout_E[44]),
    .I1(Dout_D[44]),
    .I2(_140_[0]),
    .O(_067_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _188_ (
    .I0(Dout_E[45]),
    .I1(Dout_D[45]),
    .I2(_140_[0]),
    .O(_068_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _189_ (
    .I0(Dout_E[46]),
    .I1(Dout_D[46]),
    .I2(_140_[0]),
    .O(_069_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _190_ (
    .I0(Dout_E[47]),
    .I1(Dout_D[47]),
    .I2(_140_[0]),
    .O(_070_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _191_ (
    .I0(Dout_E[48]),
    .I1(Dout_D[48]),
    .I2(_140_[0]),
    .O(_071_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _192_ (
    .I0(Dout_E[49]),
    .I1(Dout_D[49]),
    .I2(_140_[0]),
    .O(_072_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _193_ (
    .I0(Dout_E[50]),
    .I1(Dout_D[50]),
    .I2(_140_[0]),
    .O(_074_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _194_ (
    .I0(Dout_E[51]),
    .I1(Dout_D[51]),
    .I2(_140_[0]),
    .O(_075_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _195_ (
    .I0(Dout_E[52]),
    .I1(Dout_D[52]),
    .I2(_140_[0]),
    .O(_076_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _196_ (
    .I0(Dout_E[53]),
    .I1(Dout_D[53]),
    .I2(_140_[0]),
    .O(_077_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _197_ (
    .I0(Dout_E[54]),
    .I1(Dout_D[54]),
    .I2(_140_[0]),
    .O(_078_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _198_ (
    .I0(Dout_E[55]),
    .I1(Dout_D[55]),
    .I2(_140_[0]),
    .O(_079_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _199_ (
    .I0(Dout_E[56]),
    .I1(Dout_D[56]),
    .I2(_140_[0]),
    .O(_080_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _200_ (
    .I0(Dout_E[57]),
    .I1(Dout_D[57]),
    .I2(_140_[0]),
    .O(_081_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _201_ (
    .I0(Dout_E[58]),
    .I1(Dout_D[58]),
    .I2(_140_[0]),
    .O(_082_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _202_ (
    .I0(Dout_E[59]),
    .I1(Dout_D[59]),
    .I2(_140_[0]),
    .O(_083_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _203_ (
    .I0(Dout_E[60]),
    .I1(Dout_D[60]),
    .I2(_140_[0]),
    .O(_085_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _204_ (
    .I0(Dout_E[61]),
    .I1(Dout_D[61]),
    .I2(_140_[0]),
    .O(_086_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _205_ (
    .I0(Dout_E[62]),
    .I1(Dout_D[62]),
    .I2(_140_[0]),
    .O(_087_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _206_ (
    .I0(Dout_E[63]),
    .I1(Dout_D[63]),
    .I2(_140_[0]),
    .O(_088_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _207_ (
    .I0(Dout_E[64]),
    .I1(Dout_D[64]),
    .I2(_140_[0]),
    .O(_089_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _208_ (
    .I0(Dout_E[65]),
    .I1(Dout_D[65]),
    .I2(_140_[0]),
    .O(_090_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _209_ (
    .I0(Dout_E[66]),
    .I1(Dout_D[66]),
    .I2(_140_[0]),
    .O(_091_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _210_ (
    .I0(Dout_E[67]),
    .I1(Dout_D[67]),
    .I2(_140_[0]),
    .O(_092_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _211_ (
    .I0(Dout_E[68]),
    .I1(Dout_D[68]),
    .I2(_140_[0]),
    .O(_093_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _212_ (
    .I0(Dout_E[69]),
    .I1(Dout_D[69]),
    .I2(_140_[0]),
    .O(_094_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _213_ (
    .I0(Dout_E[70]),
    .I1(Dout_D[70]),
    .I2(_140_[0]),
    .O(_096_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _214_ (
    .I0(Dout_E[71]),
    .I1(Dout_D[71]),
    .I2(_140_[0]),
    .O(_097_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _215_ (
    .I0(Dout_E[72]),
    .I1(Dout_D[72]),
    .I2(_140_[0]),
    .O(_098_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _216_ (
    .I0(Dout_E[73]),
    .I1(Dout_D[73]),
    .I2(_140_[0]),
    .O(_099_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _217_ (
    .I0(Dout_E[74]),
    .I1(Dout_D[74]),
    .I2(_140_[0]),
    .O(_100_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _218_ (
    .I0(Dout_E[75]),
    .I1(Dout_D[75]),
    .I2(_140_[0]),
    .O(_101_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _219_ (
    .I0(Dout_E[76]),
    .I1(Dout_D[76]),
    .I2(_140_[0]),
    .O(_102_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _220_ (
    .I0(Dout_E[77]),
    .I1(Dout_D[77]),
    .I2(_140_[0]),
    .O(_103_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _221_ (
    .I0(Dout_E[78]),
    .I1(Dout_D[78]),
    .I2(_140_[0]),
    .O(_104_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _222_ (
    .I0(Dout_E[79]),
    .I1(Dout_D[79]),
    .I2(_140_[0]),
    .O(_105_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _223_ (
    .I0(Dout_E[80]),
    .I1(Dout_D[80]),
    .I2(_140_[0]),
    .O(_107_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _224_ (
    .I0(Dout_E[81]),
    .I1(Dout_D[81]),
    .I2(_140_[0]),
    .O(_108_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _225_ (
    .I0(Dout_E[82]),
    .I1(Dout_D[82]),
    .I2(_140_[0]),
    .O(_109_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _226_ (
    .I0(Dout_E[83]),
    .I1(Dout_D[83]),
    .I2(_140_[0]),
    .O(_110_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _227_ (
    .I0(Dout_E[84]),
    .I1(Dout_D[84]),
    .I2(_140_[0]),
    .O(_111_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _228_ (
    .I0(Dout_E[85]),
    .I1(Dout_D[85]),
    .I2(_140_[0]),
    .O(_112_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _229_ (
    .I0(Dout_E[86]),
    .I1(Dout_D[86]),
    .I2(_140_[0]),
    .O(_113_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _230_ (
    .I0(Dout_E[87]),
    .I1(Dout_D[87]),
    .I2(_140_[0]),
    .O(_114_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _231_ (
    .I0(Dout_E[88]),
    .I1(Dout_D[88]),
    .I2(_140_[0]),
    .O(_115_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _232_ (
    .I0(Dout_E[89]),
    .I1(Dout_D[89]),
    .I2(_140_[0]),
    .O(_116_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _233_ (
    .I0(Dout_E[90]),
    .I1(Dout_D[90]),
    .I2(_140_[0]),
    .O(_118_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _234_ (
    .I0(Dout_E[91]),
    .I1(Dout_D[91]),
    .I2(_140_[0]),
    .O(_119_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _235_ (
    .I0(Dout_E[92]),
    .I1(Dout_D[92]),
    .I2(_140_[0]),
    .O(_120_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _236_ (
    .I0(Dout_E[93]),
    .I1(Dout_D[93]),
    .I2(_140_[0]),
    .O(_121_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _237_ (
    .I0(Dout_E[94]),
    .I1(Dout_D[94]),
    .I2(_140_[0]),
    .O(_122_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _238_ (
    .I0(Dout_E[95]),
    .I1(Dout_D[95]),
    .I2(_140_[0]),
    .O(_123_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _239_ (
    .I0(Dout_E[96]),
    .I1(Dout_D[96]),
    .I2(_140_[0]),
    .O(_124_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _240_ (
    .I0(Dout_E[97]),
    .I1(Dout_D[97]),
    .I2(_140_[0]),
    .O(_125_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _241_ (
    .I0(Dout_E[98]),
    .I1(Dout_D[98]),
    .I2(_140_[0]),
    .O(_126_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _242_ (
    .I0(Dout_E[99]),
    .I1(Dout_D[99]),
    .I2(_140_[0]),
    .O(_127_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _243_ (
    .I0(Dout_E[100]),
    .I1(Dout_D[100]),
    .I2(_140_[0]),
    .O(_002_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _244_ (
    .I0(Dout_E[101]),
    .I1(Dout_D[101]),
    .I2(_140_[0]),
    .O(_003_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _245_ (
    .I0(Dout_E[102]),
    .I1(Dout_D[102]),
    .I2(_140_[0]),
    .O(_004_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _246_ (
    .I0(Dout_E[103]),
    .I1(Dout_D[103]),
    .I2(_140_[0]),
    .O(_005_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _247_ (
    .I0(Dout_E[104]),
    .I1(Dout_D[104]),
    .I2(_140_[0]),
    .O(_006_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _248_ (
    .I0(Dout_E[105]),
    .I1(Dout_D[105]),
    .I2(_140_[0]),
    .O(_007_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _249_ (
    .I0(Dout_E[106]),
    .I1(Dout_D[106]),
    .I2(_140_[0]),
    .O(_008_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _250_ (
    .I0(Dout_E[107]),
    .I1(Dout_D[107]),
    .I2(_140_[0]),
    .O(_009_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _251_ (
    .I0(Dout_E[108]),
    .I1(Dout_D[108]),
    .I2(_140_[0]),
    .O(_010_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _252_ (
    .I0(Dout_E[109]),
    .I1(Dout_D[109]),
    .I2(_140_[0]),
    .O(_011_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _253_ (
    .I0(Dout_E[110]),
    .I1(Dout_D[110]),
    .I2(_140_[0]),
    .O(_013_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _254_ (
    .I0(Dout_E[111]),
    .I1(Dout_D[111]),
    .I2(_140_[0]),
    .O(_014_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _255_ (
    .I0(Dout_E[112]),
    .I1(Dout_D[112]),
    .I2(_140_[0]),
    .O(_015_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _256_ (
    .I0(Dout_E[113]),
    .I1(Dout_D[113]),
    .I2(_140_[0]),
    .O(_016_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _257_ (
    .I0(Dout_E[114]),
    .I1(Dout_D[114]),
    .I2(_140_[0]),
    .O(_017_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _258_ (
    .I0(Dout_E[115]),
    .I1(Dout_D[115]),
    .I2(_140_[0]),
    .O(_018_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _259_ (
    .I0(Dout_E[116]),
    .I1(Dout_D[116]),
    .I2(_140_[0]),
    .O(_019_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _260_ (
    .I0(Dout_E[117]),
    .I1(Dout_D[117]),
    .I2(_140_[0]),
    .O(_020_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _261_ (
    .I0(Dout_E[118]),
    .I1(Dout_D[118]),
    .I2(_140_[0]),
    .O(_021_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _262_ (
    .I0(Dout_E[119]),
    .I1(Dout_D[119]),
    .I2(_140_[0]),
    .O(_022_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _263_ (
    .I0(Dout_E[120]),
    .I1(Dout_D[120]),
    .I2(_140_[0]),
    .O(_024_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _264_ (
    .I0(Dout_E[121]),
    .I1(Dout_D[121]),
    .I2(_140_[0]),
    .O(_025_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _265_ (
    .I0(Dout_E[122]),
    .I1(Dout_D[122]),
    .I2(_140_[0]),
    .O(_026_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _266_ (
    .I0(Dout_E[123]),
    .I1(Dout_D[123]),
    .I2(_140_[0]),
    .O(_027_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _267_ (
    .I0(Dout_E[124]),
    .I1(Dout_D[124]),
    .I2(_140_[0]),
    .O(_028_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _268_ (
    .I0(Dout_E[125]),
    .I1(Dout_D[125]),
    .I2(_140_[0]),
    .O(_029_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _269_ (
    .I0(Dout_E[126]),
    .I1(Dout_D[126]),
    .I2(_140_[0]),
    .O(_030_)
  );
LUT3  #(
    .INIT(8'hca)
  ) _270_ (
    .I0(Dout_E[127]),
    .I1(Dout_D[127]),
    .I2(_140_[0]),
    .O(_031_)
  );
LUT2  #(
    .INIT(4'h4)
  ) _271_ (
    .I0(_140_[0]),
    .I1(_140_[1]),
    .O(EN_E)
  );
LUT2  #(
    .INIT(4'h8)
  ) _272_ (
    .I0(_140_[0]),
    .I1(_140_[1]),
    .O(EN_D)
  );
LUT2  #(
    .INIT(4'he)
  ) _273_ (
    .I0(BSY_E),
    .I1(BSY_D),
    .O(_000_)
  );
BUFG  _274_ (
    .I(_131_),
    .O(_134_)
  );
FDRE  #(
    .INIT(1'hx)
  ) _275_ (
    .C(_134_),
    .CE(1'h1),
    .D(_133_),
    .Q(Dvld_reg),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _276_ (
    .C(_134_),
    .CE(1'h1),
    .D(_132_),
    .Q(Kvld_reg),
    .R(1'h0)
  );
LUT6  #(
    .INIT(64'ha8a80808a808a808)
  ) _277_ (
    .I0(_139_),
    .I1(Kvld_reg),
    .I2(_140_[1]),
    .I3(Kvld_E),
    .I4(Kvld_D),
    .I5(_140_[0]),
    .O(_132_)
  );
LUT6  #(
    .INIT(64'ha8a80808a808a808)
  ) _278_ (
    .I0(_139_),
    .I1(Dvld_reg),
    .I2(_140_[1]),
    .I3(Dvld_E),
    .I4(Dvld_D),
    .I5(_140_[0]),
    .O(_133_)
  );
OBUF  _279_ (
    .I(_000_),
    .O(BSY)
  );
IBUF  _280_ (
    .I(CLK),
    .O(_131_)
  );
IBUF  _281_ (
    .I(Din[0]),
    .O(_135_[0])
  );
IBUF  _282_ (
    .I(Din[1]),
    .O(_135_[1])
  );
IBUF  _283_ (
    .I(Din[10]),
    .O(_135_[10])
  );
IBUF  _284_ (
    .I(Din[100]),
    .O(_135_[100])
  );
IBUF  _285_ (
    .I(Din[101]),
    .O(_135_[101])
  );
IBUF  _286_ (
    .I(Din[102]),
    .O(_135_[102])
  );
IBUF  _287_ (
    .I(Din[103]),
    .O(_135_[103])
  );
IBUF  _288_ (
    .I(Din[104]),
    .O(_135_[104])
  );
IBUF  _289_ (
    .I(Din[105]),
    .O(_135_[105])
  );
IBUF  _290_ (
    .I(Din[106]),
    .O(_135_[106])
  );
IBUF  _291_ (
    .I(Din[107]),
    .O(_135_[107])
  );
IBUF  _292_ (
    .I(Din[108]),
    .O(_135_[108])
  );
IBUF  _293_ (
    .I(Din[109]),
    .O(_135_[109])
  );
IBUF  _294_ (
    .I(Din[11]),
    .O(_135_[11])
  );
IBUF  _295_ (
    .I(Din[110]),
    .O(_135_[110])
  );
IBUF  _296_ (
    .I(Din[111]),
    .O(_135_[111])
  );
IBUF  _297_ (
    .I(Din[112]),
    .O(_135_[112])
  );
IBUF  _298_ (
    .I(Din[113]),
    .O(_135_[113])
  );
IBUF  _299_ (
    .I(Din[114]),
    .O(_135_[114])
  );
IBUF  _300_ (
    .I(Din[115]),
    .O(_135_[115])
  );
IBUF  _301_ (
    .I(Din[116]),
    .O(_135_[116])
  );
IBUF  _302_ (
    .I(Din[117]),
    .O(_135_[117])
  );
IBUF  _303_ (
    .I(Din[118]),
    .O(_135_[118])
  );
IBUF  _304_ (
    .I(Din[119]),
    .O(_135_[119])
  );
IBUF  _305_ (
    .I(Din[12]),
    .O(_135_[12])
  );
IBUF  _306_ (
    .I(Din[120]),
    .O(_135_[120])
  );
IBUF  _307_ (
    .I(Din[121]),
    .O(_135_[121])
  );
IBUF  _308_ (
    .I(Din[122]),
    .O(_135_[122])
  );
IBUF  _309_ (
    .I(Din[123]),
    .O(_135_[123])
  );
IBUF  _310_ (
    .I(Din[124]),
    .O(_135_[124])
  );
IBUF  _311_ (
    .I(Din[125]),
    .O(_135_[125])
  );
IBUF  _312_ (
    .I(Din[126]),
    .O(_135_[126])
  );
IBUF  _313_ (
    .I(Din[127]),
    .O(_135_[127])
  );
IBUF  _314_ (
    .I(Din[13]),
    .O(_135_[13])
  );
IBUF  _315_ (
    .I(Din[14]),
    .O(_135_[14])
  );
IBUF  _316_ (
    .I(Din[15]),
    .O(_135_[15])
  );
IBUF  _317_ (
    .I(Din[16]),
    .O(_135_[16])
  );
IBUF  _318_ (
    .I(Din[17]),
    .O(_135_[17])
  );
IBUF  _319_ (
    .I(Din[18]),
    .O(_135_[18])
  );
IBUF  _320_ (
    .I(Din[19]),
    .O(_135_[19])
  );
IBUF  _321_ (
    .I(Din[2]),
    .O(_135_[2])
  );
IBUF  _322_ (
    .I(Din[20]),
    .O(_135_[20])
  );
IBUF  _323_ (
    .I(Din[21]),
    .O(_135_[21])
  );
IBUF  _324_ (
    .I(Din[22]),
    .O(_135_[22])
  );
IBUF  _325_ (
    .I(Din[23]),
    .O(_135_[23])
  );
IBUF  _326_ (
    .I(Din[24]),
    .O(_135_[24])
  );
IBUF  _327_ (
    .I(Din[25]),
    .O(_135_[25])
  );
IBUF  _328_ (
    .I(Din[26]),
    .O(_135_[26])
  );
IBUF  _329_ (
    .I(Din[27]),
    .O(_135_[27])
  );
IBUF  _330_ (
    .I(Din[28]),
    .O(_135_[28])
  );
IBUF  _331_ (
    .I(Din[29]),
    .O(_135_[29])
  );
IBUF  _332_ (
    .I(Din[3]),
    .O(_135_[3])
  );
IBUF  _333_ (
    .I(Din[30]),
    .O(_135_[30])
  );
IBUF  _334_ (
    .I(Din[31]),
    .O(_135_[31])
  );
IBUF  _335_ (
    .I(Din[32]),
    .O(_135_[32])
  );
IBUF  _336_ (
    .I(Din[33]),
    .O(_135_[33])
  );
IBUF  _337_ (
    .I(Din[34]),
    .O(_135_[34])
  );
IBUF  _338_ (
    .I(Din[35]),
    .O(_135_[35])
  );
IBUF  _339_ (
    .I(Din[36]),
    .O(_135_[36])
  );
IBUF  _340_ (
    .I(Din[37]),
    .O(_135_[37])
  );
IBUF  _341_ (
    .I(Din[38]),
    .O(_135_[38])
  );
IBUF  _342_ (
    .I(Din[39]),
    .O(_135_[39])
  );
IBUF  _343_ (
    .I(Din[4]),
    .O(_135_[4])
  );
IBUF  _344_ (
    .I(Din[40]),
    .O(_135_[40])
  );
IBUF  _345_ (
    .I(Din[41]),
    .O(_135_[41])
  );
IBUF  _346_ (
    .I(Din[42]),
    .O(_135_[42])
  );
IBUF  _347_ (
    .I(Din[43]),
    .O(_135_[43])
  );
IBUF  _348_ (
    .I(Din[44]),
    .O(_135_[44])
  );
IBUF  _349_ (
    .I(Din[45]),
    .O(_135_[45])
  );
IBUF  _350_ (
    .I(Din[46]),
    .O(_135_[46])
  );
IBUF  _351_ (
    .I(Din[47]),
    .O(_135_[47])
  );
IBUF  _352_ (
    .I(Din[48]),
    .O(_135_[48])
  );
IBUF  _353_ (
    .I(Din[49]),
    .O(_135_[49])
  );
IBUF  _354_ (
    .I(Din[5]),
    .O(_135_[5])
  );
IBUF  _355_ (
    .I(Din[50]),
    .O(_135_[50])
  );
IBUF  _356_ (
    .I(Din[51]),
    .O(_135_[51])
  );
IBUF  _357_ (
    .I(Din[52]),
    .O(_135_[52])
  );
IBUF  _358_ (
    .I(Din[53]),
    .O(_135_[53])
  );
IBUF  _359_ (
    .I(Din[54]),
    .O(_135_[54])
  );
IBUF  _360_ (
    .I(Din[55]),
    .O(_135_[55])
  );
IBUF  _361_ (
    .I(Din[56]),
    .O(_135_[56])
  );
IBUF  _362_ (
    .I(Din[57]),
    .O(_135_[57])
  );
IBUF  _363_ (
    .I(Din[58]),
    .O(_135_[58])
  );
IBUF  _364_ (
    .I(Din[59]),
    .O(_135_[59])
  );
IBUF  _365_ (
    .I(Din[6]),
    .O(_135_[6])
  );
IBUF  _366_ (
    .I(Din[60]),
    .O(_135_[60])
  );
IBUF  _367_ (
    .I(Din[61]),
    .O(_135_[61])
  );
IBUF  _368_ (
    .I(Din[62]),
    .O(_135_[62])
  );
IBUF  _369_ (
    .I(Din[63]),
    .O(_135_[63])
  );
IBUF  _370_ (
    .I(Din[64]),
    .O(_135_[64])
  );
IBUF  _371_ (
    .I(Din[65]),
    .O(_135_[65])
  );
IBUF  _372_ (
    .I(Din[66]),
    .O(_135_[66])
  );
IBUF  _373_ (
    .I(Din[67]),
    .O(_135_[67])
  );
IBUF  _374_ (
    .I(Din[68]),
    .O(_135_[68])
  );
IBUF  _375_ (
    .I(Din[69]),
    .O(_135_[69])
  );
IBUF  _376_ (
    .I(Din[7]),
    .O(_135_[7])
  );
IBUF  _377_ (
    .I(Din[70]),
    .O(_135_[70])
  );
IBUF  _378_ (
    .I(Din[71]),
    .O(_135_[71])
  );
IBUF  _379_ (
    .I(Din[72]),
    .O(_135_[72])
  );
IBUF  _380_ (
    .I(Din[73]),
    .O(_135_[73])
  );
IBUF  _381_ (
    .I(Din[74]),
    .O(_135_[74])
  );
IBUF  _382_ (
    .I(Din[75]),
    .O(_135_[75])
  );
IBUF  _383_ (
    .I(Din[76]),
    .O(_135_[76])
  );
IBUF  _384_ (
    .I(Din[77]),
    .O(_135_[77])
  );
IBUF  _385_ (
    .I(Din[78]),
    .O(_135_[78])
  );
IBUF  _386_ (
    .I(Din[79]),
    .O(_135_[79])
  );
IBUF  _387_ (
    .I(Din[8]),
    .O(_135_[8])
  );
IBUF  _388_ (
    .I(Din[80]),
    .O(_135_[80])
  );
IBUF  _389_ (
    .I(Din[81]),
    .O(_135_[81])
  );
IBUF  _390_ (
    .I(Din[82]),
    .O(_135_[82])
  );
IBUF  _391_ (
    .I(Din[83]),
    .O(_135_[83])
  );
IBUF  _392_ (
    .I(Din[84]),
    .O(_135_[84])
  );
IBUF  _393_ (
    .I(Din[85]),
    .O(_135_[85])
  );
IBUF  _394_ (
    .I(Din[86]),
    .O(_135_[86])
  );
IBUF  _395_ (
    .I(Din[87]),
    .O(_135_[87])
  );
IBUF  _396_ (
    .I(Din[88]),
    .O(_135_[88])
  );
IBUF  _397_ (
    .I(Din[89]),
    .O(_135_[89])
  );
IBUF  _398_ (
    .I(Din[9]),
    .O(_135_[9])
  );
IBUF  _399_ (
    .I(Din[90]),
    .O(_135_[90])
  );
IBUF  _400_ (
    .I(Din[91]),
    .O(_135_[91])
  );
IBUF  _401_ (
    .I(Din[92]),
    .O(_135_[92])
  );
IBUF  _402_ (
    .I(Din[93]),
    .O(_135_[93])
  );
IBUF  _403_ (
    .I(Din[94]),
    .O(_135_[94])
  );
IBUF  _404_ (
    .I(Din[95]),
    .O(_135_[95])
  );
IBUF  _405_ (
    .I(Din[96]),
    .O(_135_[96])
  );
IBUF  _406_ (
    .I(Din[97]),
    .O(_135_[97])
  );
IBUF  _407_ (
    .I(Din[98]),
    .O(_135_[98])
  );
IBUF  _408_ (
    .I(Din[99]),
    .O(_135_[99])
  );
OBUF  _409_ (
    .I(_001_),
    .O(Dout[0])
  );
OBUF  _410_ (
    .I(_040_),
    .O(Dout[1])
  );
OBUF  _411_ (
    .I(_012_),
    .O(Dout[10])
  );
OBUF  _412_ (
    .I(_002_),
    .O(Dout[100])
  );
OBUF  _413_ (
    .I(_003_),
    .O(Dout[101])
  );
OBUF  _414_ (
    .I(_004_),
    .O(Dout[102])
  );
OBUF  _415_ (
    .I(_005_),
    .O(Dout[103])
  );
OBUF  _416_ (
    .I(_006_),
    .O(Dout[104])
  );
OBUF  _417_ (
    .I(_007_),
    .O(Dout[105])
  );
OBUF  _418_ (
    .I(_008_),
    .O(Dout[106])
  );
OBUF  _419_ (
    .I(_009_),
    .O(Dout[107])
  );
OBUF  _420_ (
    .I(_010_),
    .O(Dout[108])
  );
OBUF  _421_ (
    .I(_011_),
    .O(Dout[109])
  );
OBUF  _422_ (
    .I(_023_),
    .O(Dout[11])
  );
OBUF  _423_ (
    .I(_013_),
    .O(Dout[110])
  );
OBUF  _424_ (
    .I(_014_),
    .O(Dout[111])
  );
OBUF  _425_ (
    .I(_015_),
    .O(Dout[112])
  );
OBUF  _426_ (
    .I(_016_),
    .O(Dout[113])
  );
OBUF  _427_ (
    .I(_017_),
    .O(Dout[114])
  );
OBUF  _428_ (
    .I(_018_),
    .O(Dout[115])
  );
OBUF  _429_ (
    .I(_019_),
    .O(Dout[116])
  );
OBUF  _430_ (
    .I(_020_),
    .O(Dout[117])
  );
OBUF  _431_ (
    .I(_021_),
    .O(Dout[118])
  );
OBUF  _432_ (
    .I(_022_),
    .O(Dout[119])
  );
OBUF  _433_ (
    .I(_032_),
    .O(Dout[12])
  );
OBUF  _434_ (
    .I(_024_),
    .O(Dout[120])
  );
OBUF  _435_ (
    .I(_025_),
    .O(Dout[121])
  );
OBUF  _436_ (
    .I(_026_),
    .O(Dout[122])
  );
OBUF  _437_ (
    .I(_027_),
    .O(Dout[123])
  );
OBUF  _438_ (
    .I(_028_),
    .O(Dout[124])
  );
OBUF  _439_ (
    .I(_029_),
    .O(Dout[125])
  );
OBUF  _440_ (
    .I(_030_),
    .O(Dout[126])
  );
OBUF  _441_ (
    .I(_031_),
    .O(Dout[127])
  );
OBUF  _442_ (
    .I(_033_),
    .O(Dout[13])
  );
OBUF  _443_ (
    .I(_034_),
    .O(Dout[14])
  );
OBUF  _444_ (
    .I(_035_),
    .O(Dout[15])
  );
OBUF  _445_ (
    .I(_036_),
    .O(Dout[16])
  );
OBUF  _446_ (
    .I(_037_),
    .O(Dout[17])
  );
OBUF  _447_ (
    .I(_038_),
    .O(Dout[18])
  );
OBUF  _448_ (
    .I(_039_),
    .O(Dout[19])
  );
OBUF  _449_ (
    .I(_051_),
    .O(Dout[2])
  );
OBUF  _450_ (
    .I(_041_),
    .O(Dout[20])
  );
OBUF  _451_ (
    .I(_042_),
    .O(Dout[21])
  );
OBUF  _452_ (
    .I(_043_),
    .O(Dout[22])
  );
OBUF  _453_ (
    .I(_044_),
    .O(Dout[23])
  );
OBUF  _454_ (
    .I(_045_),
    .O(Dout[24])
  );
OBUF  _455_ (
    .I(_046_),
    .O(Dout[25])
  );
OBUF  _456_ (
    .I(_047_),
    .O(Dout[26])
  );
OBUF  _457_ (
    .I(_048_),
    .O(Dout[27])
  );
OBUF  _458_ (
    .I(_049_),
    .O(Dout[28])
  );
OBUF  _459_ (
    .I(_050_),
    .O(Dout[29])
  );
OBUF  _460_ (
    .I(_062_),
    .O(Dout[3])
  );
OBUF  _461_ (
    .I(_052_),
    .O(Dout[30])
  );
OBUF  _462_ (
    .I(_053_),
    .O(Dout[31])
  );
OBUF  _463_ (
    .I(_054_),
    .O(Dout[32])
  );
OBUF  _464_ (
    .I(_055_),
    .O(Dout[33])
  );
OBUF  _465_ (
    .I(_056_),
    .O(Dout[34])
  );
OBUF  _466_ (
    .I(_057_),
    .O(Dout[35])
  );
OBUF  _467_ (
    .I(_058_),
    .O(Dout[36])
  );
OBUF  _468_ (
    .I(_059_),
    .O(Dout[37])
  );
OBUF  _469_ (
    .I(_060_),
    .O(Dout[38])
  );
OBUF  _470_ (
    .I(_061_),
    .O(Dout[39])
  );
OBUF  _471_ (
    .I(_073_),
    .O(Dout[4])
  );
OBUF  _472_ (
    .I(_063_),
    .O(Dout[40])
  );
OBUF  _473_ (
    .I(_064_),
    .O(Dout[41])
  );
OBUF  _474_ (
    .I(_065_),
    .O(Dout[42])
  );
OBUF  _475_ (
    .I(_066_),
    .O(Dout[43])
  );
OBUF  _476_ (
    .I(_067_),
    .O(Dout[44])
  );
OBUF  _477_ (
    .I(_068_),
    .O(Dout[45])
  );
OBUF  _478_ (
    .I(_069_),
    .O(Dout[46])
  );
OBUF  _479_ (
    .I(_070_),
    .O(Dout[47])
  );
OBUF  _480_ (
    .I(_071_),
    .O(Dout[48])
  );
OBUF  _481_ (
    .I(_072_),
    .O(Dout[49])
  );
OBUF  _482_ (
    .I(_084_),
    .O(Dout[5])
  );
OBUF  _483_ (
    .I(_074_),
    .O(Dout[50])
  );
OBUF  _484_ (
    .I(_075_),
    .O(Dout[51])
  );
OBUF  _485_ (
    .I(_076_),
    .O(Dout[52])
  );
OBUF  _486_ (
    .I(_077_),
    .O(Dout[53])
  );
OBUF  _487_ (
    .I(_078_),
    .O(Dout[54])
  );
OBUF  _488_ (
    .I(_079_),
    .O(Dout[55])
  );
OBUF  _489_ (
    .I(_080_),
    .O(Dout[56])
  );
OBUF  _490_ (
    .I(_081_),
    .O(Dout[57])
  );
OBUF  _491_ (
    .I(_082_),
    .O(Dout[58])
  );
OBUF  _492_ (
    .I(_083_),
    .O(Dout[59])
  );
OBUF  _493_ (
    .I(_095_),
    .O(Dout[6])
  );
OBUF  _494_ (
    .I(_085_),
    .O(Dout[60])
  );
OBUF  _495_ (
    .I(_086_),
    .O(Dout[61])
  );
OBUF  _496_ (
    .I(_087_),
    .O(Dout[62])
  );
OBUF  _497_ (
    .I(_088_),
    .O(Dout[63])
  );
OBUF  _498_ (
    .I(_089_),
    .O(Dout[64])
  );
OBUF  _499_ (
    .I(_090_),
    .O(Dout[65])
  );
OBUF  _500_ (
    .I(_091_),
    .O(Dout[66])
  );
OBUF  _501_ (
    .I(_092_),
    .O(Dout[67])
  );
OBUF  _502_ (
    .I(_093_),
    .O(Dout[68])
  );
OBUF  _503_ (
    .I(_094_),
    .O(Dout[69])
  );
OBUF  _504_ (
    .I(_106_),
    .O(Dout[7])
  );
OBUF  _505_ (
    .I(_096_),
    .O(Dout[70])
  );
OBUF  _506_ (
    .I(_097_),
    .O(Dout[71])
  );
OBUF  _507_ (
    .I(_098_),
    .O(Dout[72])
  );
OBUF  _508_ (
    .I(_099_),
    .O(Dout[73])
  );
OBUF  _509_ (
    .I(_100_),
    .O(Dout[74])
  );
OBUF  _510_ (
    .I(_101_),
    .O(Dout[75])
  );
OBUF  _511_ (
    .I(_102_),
    .O(Dout[76])
  );
OBUF  _512_ (
    .I(_103_),
    .O(Dout[77])
  );
OBUF  _513_ (
    .I(_104_),
    .O(Dout[78])
  );
OBUF  _514_ (
    .I(_105_),
    .O(Dout[79])
  );
OBUF  _515_ (
    .I(_117_),
    .O(Dout[8])
  );
OBUF  _516_ (
    .I(_107_),
    .O(Dout[80])
  );
OBUF  _517_ (
    .I(_108_),
    .O(Dout[81])
  );
OBUF  _518_ (
    .I(_109_),
    .O(Dout[82])
  );
OBUF  _519_ (
    .I(_110_),
    .O(Dout[83])
  );
OBUF  _520_ (
    .I(_111_),
    .O(Dout[84])
  );
OBUF  _521_ (
    .I(_112_),
    .O(Dout[85])
  );
OBUF  _522_ (
    .I(_113_),
    .O(Dout[86])
  );
OBUF  _523_ (
    .I(_114_),
    .O(Dout[87])
  );
OBUF  _524_ (
    .I(_115_),
    .O(Dout[88])
  );
OBUF  _525_ (
    .I(_116_),
    .O(Dout[89])
  );
OBUF  _526_ (
    .I(_128_),
    .O(Dout[9])
  );
OBUF  _527_ (
    .I(_118_),
    .O(Dout[90])
  );
OBUF  _528_ (
    .I(_119_),
    .O(Dout[91])
  );
OBUF  _529_ (
    .I(_120_),
    .O(Dout[92])
  );
OBUF  _530_ (
    .I(_121_),
    .O(Dout[93])
  );
OBUF  _531_ (
    .I(_122_),
    .O(Dout[94])
  );
OBUF  _532_ (
    .I(_123_),
    .O(Dout[95])
  );
OBUF  _533_ (
    .I(_124_),
    .O(Dout[96])
  );
OBUF  _534_ (
    .I(_125_),
    .O(Dout[97])
  );
OBUF  _535_ (
    .I(_126_),
    .O(Dout[98])
  );
OBUF  _536_ (
    .I(_127_),
    .O(Dout[99])
  );
IBUF  _537_ (
    .I(Drdy),
    .O(_136_)
  );
OBUF  _538_ (
    .I(_129_),
    .O(Dvld)
  );
IBUF  _539_ (
    .I(EN),
    .O(_140_[1])
  );
IBUF  _540_ (
    .I(EncDec),
    .O(_140_[0])
  );
IBUF  _541_ (
    .I(Kin[0]),
    .O(_137_[0])
  );
IBUF  _542_ (
    .I(Kin[1]),
    .O(_137_[1])
  );
IBUF  _543_ (
    .I(Kin[10]),
    .O(_137_[10])
  );
IBUF  _544_ (
    .I(Kin[100]),
    .O(_137_[100])
  );
IBUF  _545_ (
    .I(Kin[101]),
    .O(_137_[101])
  );
IBUF  _546_ (
    .I(Kin[102]),
    .O(_137_[102])
  );
IBUF  _547_ (
    .I(Kin[103]),
    .O(_137_[103])
  );
IBUF  _548_ (
    .I(Kin[104]),
    .O(_137_[104])
  );
IBUF  _549_ (
    .I(Kin[105]),
    .O(_137_[105])
  );
IBUF  _550_ (
    .I(Kin[106]),
    .O(_137_[106])
  );
IBUF  _551_ (
    .I(Kin[107]),
    .O(_137_[107])
  );
IBUF  _552_ (
    .I(Kin[108]),
    .O(_137_[108])
  );
IBUF  _553_ (
    .I(Kin[109]),
    .O(_137_[109])
  );
IBUF  _554_ (
    .I(Kin[11]),
    .O(_137_[11])
  );
IBUF  _555_ (
    .I(Kin[110]),
    .O(_137_[110])
  );
IBUF  _556_ (
    .I(Kin[111]),
    .O(_137_[111])
  );
IBUF  _557_ (
    .I(Kin[112]),
    .O(_137_[112])
  );
IBUF  _558_ (
    .I(Kin[113]),
    .O(_137_[113])
  );
IBUF  _559_ (
    .I(Kin[114]),
    .O(_137_[114])
  );
IBUF  _560_ (
    .I(Kin[115]),
    .O(_137_[115])
  );
IBUF  _561_ (
    .I(Kin[116]),
    .O(_137_[116])
  );
IBUF  _562_ (
    .I(Kin[117]),
    .O(_137_[117])
  );
IBUF  _563_ (
    .I(Kin[118]),
    .O(_137_[118])
  );
IBUF  _564_ (
    .I(Kin[119]),
    .O(_137_[119])
  );
IBUF  _565_ (
    .I(Kin[12]),
    .O(_137_[12])
  );
IBUF  _566_ (
    .I(Kin[120]),
    .O(_137_[120])
  );
IBUF  _567_ (
    .I(Kin[121]),
    .O(_137_[121])
  );
IBUF  _568_ (
    .I(Kin[122]),
    .O(_137_[122])
  );
IBUF  _569_ (
    .I(Kin[123]),
    .O(_137_[123])
  );
IBUF  _570_ (
    .I(Kin[124]),
    .O(_137_[124])
  );
IBUF  _571_ (
    .I(Kin[125]),
    .O(_137_[125])
  );
IBUF  _572_ (
    .I(Kin[126]),
    .O(_137_[126])
  );
IBUF  _573_ (
    .I(Kin[127]),
    .O(_137_[127])
  );
IBUF  _574_ (
    .I(Kin[13]),
    .O(_137_[13])
  );
IBUF  _575_ (
    .I(Kin[14]),
    .O(_137_[14])
  );
IBUF  _576_ (
    .I(Kin[15]),
    .O(_137_[15])
  );
IBUF  _577_ (
    .I(Kin[16]),
    .O(_137_[16])
  );
IBUF  _578_ (
    .I(Kin[17]),
    .O(_137_[17])
  );
IBUF  _579_ (
    .I(Kin[18]),
    .O(_137_[18])
  );
IBUF  _580_ (
    .I(Kin[19]),
    .O(_137_[19])
  );
IBUF  _581_ (
    .I(Kin[2]),
    .O(_137_[2])
  );
IBUF  _582_ (
    .I(Kin[20]),
    .O(_137_[20])
  );
IBUF  _583_ (
    .I(Kin[21]),
    .O(_137_[21])
  );
IBUF  _584_ (
    .I(Kin[22]),
    .O(_137_[22])
  );
IBUF  _585_ (
    .I(Kin[23]),
    .O(_137_[23])
  );
IBUF  _586_ (
    .I(Kin[24]),
    .O(_137_[24])
  );
IBUF  _587_ (
    .I(Kin[25]),
    .O(_137_[25])
  );
IBUF  _588_ (
    .I(Kin[26]),
    .O(_137_[26])
  );
IBUF  _589_ (
    .I(Kin[27]),
    .O(_137_[27])
  );
IBUF  _590_ (
    .I(Kin[28]),
    .O(_137_[28])
  );
IBUF  _591_ (
    .I(Kin[29]),
    .O(_137_[29])
  );
IBUF  _592_ (
    .I(Kin[3]),
    .O(_137_[3])
  );
IBUF  _593_ (
    .I(Kin[30]),
    .O(_137_[30])
  );
IBUF  _594_ (
    .I(Kin[31]),
    .O(_137_[31])
  );
IBUF  _595_ (
    .I(Kin[32]),
    .O(_137_[32])
  );
IBUF  _596_ (
    .I(Kin[33]),
    .O(_137_[33])
  );
IBUF  _597_ (
    .I(Kin[34]),
    .O(_137_[34])
  );
IBUF  _598_ (
    .I(Kin[35]),
    .O(_137_[35])
  );
IBUF  _599_ (
    .I(Kin[36]),
    .O(_137_[36])
  );
IBUF  _600_ (
    .I(Kin[37]),
    .O(_137_[37])
  );
IBUF  _601_ (
    .I(Kin[38]),
    .O(_137_[38])
  );
IBUF  _602_ (
    .I(Kin[39]),
    .O(_137_[39])
  );
IBUF  _603_ (
    .I(Kin[4]),
    .O(_137_[4])
  );
IBUF  _604_ (
    .I(Kin[40]),
    .O(_137_[40])
  );
IBUF  _605_ (
    .I(Kin[41]),
    .O(_137_[41])
  );
IBUF  _606_ (
    .I(Kin[42]),
    .O(_137_[42])
  );
IBUF  _607_ (
    .I(Kin[43]),
    .O(_137_[43])
  );
IBUF  _608_ (
    .I(Kin[44]),
    .O(_137_[44])
  );
IBUF  _609_ (
    .I(Kin[45]),
    .O(_137_[45])
  );
IBUF  _610_ (
    .I(Kin[46]),
    .O(_137_[46])
  );
IBUF  _611_ (
    .I(Kin[47]),
    .O(_137_[47])
  );
IBUF  _612_ (
    .I(Kin[48]),
    .O(_137_[48])
  );
IBUF  _613_ (
    .I(Kin[49]),
    .O(_137_[49])
  );
IBUF  _614_ (
    .I(Kin[5]),
    .O(_137_[5])
  );
IBUF  _615_ (
    .I(Kin[50]),
    .O(_137_[50])
  );
IBUF  _616_ (
    .I(Kin[51]),
    .O(_137_[51])
  );
IBUF  _617_ (
    .I(Kin[52]),
    .O(_137_[52])
  );
IBUF  _618_ (
    .I(Kin[53]),
    .O(_137_[53])
  );
IBUF  _619_ (
    .I(Kin[54]),
    .O(_137_[54])
  );
IBUF  _620_ (
    .I(Kin[55]),
    .O(_137_[55])
  );
IBUF  _621_ (
    .I(Kin[56]),
    .O(_137_[56])
  );
IBUF  _622_ (
    .I(Kin[57]),
    .O(_137_[57])
  );
IBUF  _623_ (
    .I(Kin[58]),
    .O(_137_[58])
  );
IBUF  _624_ (
    .I(Kin[59]),
    .O(_137_[59])
  );
IBUF  _625_ (
    .I(Kin[6]),
    .O(_137_[6])
  );
IBUF  _626_ (
    .I(Kin[60]),
    .O(_137_[60])
  );
IBUF  _627_ (
    .I(Kin[61]),
    .O(_137_[61])
  );
IBUF  _628_ (
    .I(Kin[62]),
    .O(_137_[62])
  );
IBUF  _629_ (
    .I(Kin[63]),
    .O(_137_[63])
  );
IBUF  _630_ (
    .I(Kin[64]),
    .O(_137_[64])
  );
IBUF  _631_ (
    .I(Kin[65]),
    .O(_137_[65])
  );
IBUF  _632_ (
    .I(Kin[66]),
    .O(_137_[66])
  );
IBUF  _633_ (
    .I(Kin[67]),
    .O(_137_[67])
  );
IBUF  _634_ (
    .I(Kin[68]),
    .O(_137_[68])
  );
IBUF  _635_ (
    .I(Kin[69]),
    .O(_137_[69])
  );
IBUF  _636_ (
    .I(Kin[7]),
    .O(_137_[7])
  );
IBUF  _637_ (
    .I(Kin[70]),
    .O(_137_[70])
  );
IBUF  _638_ (
    .I(Kin[71]),
    .O(_137_[71])
  );
IBUF  _639_ (
    .I(Kin[72]),
    .O(_137_[72])
  );
IBUF  _640_ (
    .I(Kin[73]),
    .O(_137_[73])
  );
IBUF  _641_ (
    .I(Kin[74]),
    .O(_137_[74])
  );
IBUF  _642_ (
    .I(Kin[75]),
    .O(_137_[75])
  );
IBUF  _643_ (
    .I(Kin[76]),
    .O(_137_[76])
  );
IBUF  _644_ (
    .I(Kin[77]),
    .O(_137_[77])
  );
IBUF  _645_ (
    .I(Kin[78]),
    .O(_137_[78])
  );
IBUF  _646_ (
    .I(Kin[79]),
    .O(_137_[79])
  );
IBUF  _647_ (
    .I(Kin[8]),
    .O(_137_[8])
  );
IBUF  _648_ (
    .I(Kin[80]),
    .O(_137_[80])
  );
IBUF  _649_ (
    .I(Kin[81]),
    .O(_137_[81])
  );
IBUF  _650_ (
    .I(Kin[82]),
    .O(_137_[82])
  );
IBUF  _651_ (
    .I(Kin[83]),
    .O(_137_[83])
  );
IBUF  _652_ (
    .I(Kin[84]),
    .O(_137_[84])
  );
IBUF  _653_ (
    .I(Kin[85]),
    .O(_137_[85])
  );
IBUF  _654_ (
    .I(Kin[86]),
    .O(_137_[86])
  );
IBUF  _655_ (
    .I(Kin[87]),
    .O(_137_[87])
  );
IBUF  _656_ (
    .I(Kin[88]),
    .O(_137_[88])
  );
IBUF  _657_ (
    .I(Kin[89]),
    .O(_137_[89])
  );
IBUF  _658_ (
    .I(Kin[9]),
    .O(_137_[9])
  );
IBUF  _659_ (
    .I(Kin[90]),
    .O(_137_[90])
  );
IBUF  _660_ (
    .I(Kin[91]),
    .O(_137_[91])
  );
IBUF  _661_ (
    .I(Kin[92]),
    .O(_137_[92])
  );
IBUF  _662_ (
    .I(Kin[93]),
    .O(_137_[93])
  );
IBUF  _663_ (
    .I(Kin[94]),
    .O(_137_[94])
  );
IBUF  _664_ (
    .I(Kin[95]),
    .O(_137_[95])
  );
IBUF  _665_ (
    .I(Kin[96]),
    .O(_137_[96])
  );
IBUF  _666_ (
    .I(Kin[97]),
    .O(_137_[97])
  );
IBUF  _667_ (
    .I(Kin[98]),
    .O(_137_[98])
  );
IBUF  _668_ (
    .I(Kin[99]),
    .O(_137_[99])
  );
IBUF  _669_ (
    .I(Krdy),
    .O(_138_)
  );
OBUF  _670_ (
    .I(_130_),
    .O(Kvld)
  );
IBUF  _671_ (
    .I(RSTn),
    .O(_139_)
  );
AES_Comp_DEC  AES_Comp_DEC (
    .BSY(BSY_D),
    .CLK(_134_),
    .Din(_135_),
    .Dout(Dout_D),
    .Drdy(_136_),
    .Dvld(Dvld_D),
    .EN(EN_D),
    .Kin(_137_),
    .Krdy(_138_),
    .Kvld(Kvld_D),
    .RSTn(_139_)
  );
AES_Comp_ENC  AES_Comp_ENC (
    .BSY(BSY_E),
    .CLK(_134_),
    .Din(_135_),
    .Dout(Dout_E),
    .Drdy(_136_),
    .Dvld(Dvld_E),
    .EN(EN_E),
    .Kin(_137_),
    .Krdy(_138_),
    .Kvld(Kvld_E),
    .RSTn(_139_)
  );
endmodule
