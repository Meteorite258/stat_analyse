module one_round(clk,  state_in, key, state_out);
input  clk;
wire  [31:0] k0;
wire  [31:0] k1;
wire  [31:0] k2;
wire  [31:0] k3;
input  [127:0] key;
wire  [31:0] p00;
wire  [31:0] p01;
wire  [31:0] p02;
wire  [31:0] p03;
wire  [31:0] p10;
wire  [31:0] p11;
wire  [31:0] p12;
wire  [31:0] p13;
wire  [31:0] p20;
wire  [31:0] p21;
wire  [31:0] p22;
wire  [31:0] p23;
wire  [31:0] p30;
wire  [31:0] p31;
wire  [31:0] p32;
wire  [31:0] p33;
wire  [31:0] s0;
wire  [31:0] s1;
wire  [31:0] s2;
wire  [31:0] s3;
input  [127:0] state_in;
output  [127:0] state_out;
wire  [31:0] z0;
wire  [31:0] z1;
wire  [31:0] z2;
wire  [31:0] z3;
LUT5  #(
    .INIT(32'd2523490710)
  ) _000_ (
    .I0(p00[0]),
    .I1(p11[0]),
    .I2(p22[0]),
    .I3(p33[0]),
    .I4(key[96]),
    .O(z0[0])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _001_ (
    .I0(p00[1]),
    .I1(p11[1]),
    .I2(p22[1]),
    .I3(p33[1]),
    .I4(key[97]),
    .O(z0[1])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _002_ (
    .I0(p00[2]),
    .I1(p11[2]),
    .I2(p22[2]),
    .I3(p33[2]),
    .I4(key[98]),
    .O(z0[2])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _003_ (
    .I0(p00[3]),
    .I1(p11[3]),
    .I2(p22[3]),
    .I3(p33[3]),
    .I4(key[99]),
    .O(z0[3])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _004_ (
    .I0(p00[4]),
    .I1(p11[4]),
    .I2(p22[4]),
    .I3(p33[4]),
    .I4(key[100]),
    .O(z0[4])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _005_ (
    .I0(p00[5]),
    .I1(p11[5]),
    .I2(p22[5]),
    .I3(p33[5]),
    .I4(key[101]),
    .O(z0[5])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _006_ (
    .I0(p00[6]),
    .I1(p11[6]),
    .I2(p22[6]),
    .I3(p33[6]),
    .I4(key[102]),
    .O(z0[6])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _007_ (
    .I0(p00[7]),
    .I1(p11[7]),
    .I2(p22[7]),
    .I3(p33[7]),
    .I4(key[103]),
    .O(z0[7])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _008_ (
    .I0(p00[8]),
    .I1(p11[8]),
    .I2(p22[8]),
    .I3(p33[8]),
    .I4(key[104]),
    .O(z0[8])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _009_ (
    .I0(p00[9]),
    .I1(p11[9]),
    .I2(p22[9]),
    .I3(p33[9]),
    .I4(key[105]),
    .O(z0[9])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _010_ (
    .I0(p00[10]),
    .I1(p11[10]),
    .I2(p22[10]),
    .I3(p33[10]),
    .I4(key[106]),
    .O(z0[10])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _011_ (
    .I0(p00[11]),
    .I1(p11[11]),
    .I2(p22[11]),
    .I3(p33[11]),
    .I4(key[107]),
    .O(z0[11])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _012_ (
    .I0(p00[12]),
    .I1(p11[12]),
    .I2(p22[12]),
    .I3(p33[12]),
    .I4(key[108]),
    .O(z0[12])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _013_ (
    .I0(p00[13]),
    .I1(p11[13]),
    .I2(p22[13]),
    .I3(p33[13]),
    .I4(key[109]),
    .O(z0[13])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _014_ (
    .I0(p00[14]),
    .I1(p11[14]),
    .I2(p22[14]),
    .I3(p33[14]),
    .I4(key[110]),
    .O(z0[14])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _015_ (
    .I0(p00[15]),
    .I1(p11[15]),
    .I2(p22[15]),
    .I3(p33[15]),
    .I4(key[111]),
    .O(z0[15])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _016_ (
    .I0(p00[16]),
    .I1(p11[16]),
    .I2(p22[16]),
    .I3(p33[16]),
    .I4(key[112]),
    .O(z0[16])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _017_ (
    .I0(p00[17]),
    .I1(p11[17]),
    .I2(p22[17]),
    .I3(p33[17]),
    .I4(key[113]),
    .O(z0[17])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _018_ (
    .I0(p00[18]),
    .I1(p11[18]),
    .I2(p22[18]),
    .I3(p33[18]),
    .I4(key[114]),
    .O(z0[18])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _019_ (
    .I0(p00[19]),
    .I1(p11[19]),
    .I2(p22[19]),
    .I3(p33[19]),
    .I4(key[115]),
    .O(z0[19])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _020_ (
    .I0(p00[20]),
    .I1(p11[20]),
    .I2(p22[20]),
    .I3(p33[20]),
    .I4(key[116]),
    .O(z0[20])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _021_ (
    .I0(p00[21]),
    .I1(p11[21]),
    .I2(p22[21]),
    .I3(p33[21]),
    .I4(key[117]),
    .O(z0[21])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _022_ (
    .I0(p00[22]),
    .I1(p11[22]),
    .I2(p22[22]),
    .I3(p33[22]),
    .I4(key[118]),
    .O(z0[22])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _023_ (
    .I0(p00[23]),
    .I1(p11[23]),
    .I2(p22[23]),
    .I3(p33[23]),
    .I4(key[119]),
    .O(z0[23])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _024_ (
    .I0(p00[24]),
    .I1(p11[24]),
    .I2(p22[24]),
    .I3(p33[24]),
    .I4(key[120]),
    .O(z0[24])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _025_ (
    .I0(p00[25]),
    .I1(p11[25]),
    .I2(p22[25]),
    .I3(p33[25]),
    .I4(key[121]),
    .O(z0[25])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _026_ (
    .I0(p00[26]),
    .I1(p11[26]),
    .I2(p22[26]),
    .I3(p33[26]),
    .I4(key[122]),
    .O(z0[26])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _027_ (
    .I0(p00[27]),
    .I1(p11[27]),
    .I2(p22[27]),
    .I3(p33[27]),
    .I4(key[123]),
    .O(z0[27])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _028_ (
    .I0(p00[28]),
    .I1(p11[28]),
    .I2(p22[28]),
    .I3(p33[28]),
    .I4(key[124]),
    .O(z0[28])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _029_ (
    .I0(p00[29]),
    .I1(p11[29]),
    .I2(p22[29]),
    .I3(p33[29]),
    .I4(key[125]),
    .O(z0[29])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _030_ (
    .I0(p00[30]),
    .I1(p11[30]),
    .I2(p22[30]),
    .I3(p33[30]),
    .I4(key[126]),
    .O(z0[30])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _031_ (
    .I0(p00[31]),
    .I1(p11[31]),
    .I2(p22[31]),
    .I3(p33[31]),
    .I4(key[127]),
    .O(z0[31])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _032_ (
    .I0(p03[0]),
    .I1(p10[0]),
    .I2(p21[0]),
    .I3(p32[0]),
    .I4(key[64]),
    .O(z1[0])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _033_ (
    .I0(p03[1]),
    .I1(p10[1]),
    .I2(p21[1]),
    .I3(p32[1]),
    .I4(key[65]),
    .O(z1[1])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _034_ (
    .I0(p03[2]),
    .I1(p10[2]),
    .I2(p21[2]),
    .I3(p32[2]),
    .I4(key[66]),
    .O(z1[2])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _035_ (
    .I0(p03[3]),
    .I1(p10[3]),
    .I2(p21[3]),
    .I3(p32[3]),
    .I4(key[67]),
    .O(z1[3])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _036_ (
    .I0(p03[4]),
    .I1(p10[4]),
    .I2(p21[4]),
    .I3(p32[4]),
    .I4(key[68]),
    .O(z1[4])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _037_ (
    .I0(p03[5]),
    .I1(p10[5]),
    .I2(p21[5]),
    .I3(p32[5]),
    .I4(key[69]),
    .O(z1[5])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _038_ (
    .I0(p03[6]),
    .I1(p10[6]),
    .I2(p21[6]),
    .I3(p32[6]),
    .I4(key[70]),
    .O(z1[6])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _039_ (
    .I0(p03[7]),
    .I1(p10[7]),
    .I2(p21[7]),
    .I3(p32[7]),
    .I4(key[71]),
    .O(z1[7])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _040_ (
    .I0(p03[8]),
    .I1(p10[8]),
    .I2(p21[8]),
    .I3(p32[8]),
    .I4(key[72]),
    .O(z1[8])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _041_ (
    .I0(p03[9]),
    .I1(p10[9]),
    .I2(p21[9]),
    .I3(p32[9]),
    .I4(key[73]),
    .O(z1[9])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _042_ (
    .I0(p03[10]),
    .I1(p10[10]),
    .I2(p21[10]),
    .I3(p32[10]),
    .I4(key[74]),
    .O(z1[10])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _043_ (
    .I0(p03[11]),
    .I1(p10[11]),
    .I2(p21[11]),
    .I3(p32[11]),
    .I4(key[75]),
    .O(z1[11])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _044_ (
    .I0(p03[12]),
    .I1(p10[12]),
    .I2(p21[12]),
    .I3(p32[12]),
    .I4(key[76]),
    .O(z1[12])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _045_ (
    .I0(p03[13]),
    .I1(p10[13]),
    .I2(p21[13]),
    .I3(p32[13]),
    .I4(key[77]),
    .O(z1[13])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _046_ (
    .I0(p03[14]),
    .I1(p10[14]),
    .I2(p21[14]),
    .I3(p32[14]),
    .I4(key[78]),
    .O(z1[14])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _047_ (
    .I0(p03[15]),
    .I1(p10[15]),
    .I2(p21[15]),
    .I3(p32[15]),
    .I4(key[79]),
    .O(z1[15])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _048_ (
    .I0(p03[16]),
    .I1(p10[16]),
    .I2(p21[16]),
    .I3(p32[16]),
    .I4(key[80]),
    .O(z1[16])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _049_ (
    .I0(p03[17]),
    .I1(p10[17]),
    .I2(p21[17]),
    .I3(p32[17]),
    .I4(key[81]),
    .O(z1[17])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _050_ (
    .I0(p03[18]),
    .I1(p10[18]),
    .I2(p21[18]),
    .I3(p32[18]),
    .I4(key[82]),
    .O(z1[18])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _051_ (
    .I0(p03[19]),
    .I1(p10[19]),
    .I2(p21[19]),
    .I3(p32[19]),
    .I4(key[83]),
    .O(z1[19])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _052_ (
    .I0(p03[20]),
    .I1(p10[20]),
    .I2(p21[20]),
    .I3(p32[20]),
    .I4(key[84]),
    .O(z1[20])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _053_ (
    .I0(p03[21]),
    .I1(p10[21]),
    .I2(p21[21]),
    .I3(p32[21]),
    .I4(key[85]),
    .O(z1[21])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _054_ (
    .I0(p03[22]),
    .I1(p10[22]),
    .I2(p21[22]),
    .I3(p32[22]),
    .I4(key[86]),
    .O(z1[22])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _055_ (
    .I0(p03[23]),
    .I1(p10[23]),
    .I2(p21[23]),
    .I3(p32[23]),
    .I4(key[87]),
    .O(z1[23])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _056_ (
    .I0(p03[24]),
    .I1(p10[24]),
    .I2(p21[24]),
    .I3(p32[24]),
    .I4(key[88]),
    .O(z1[24])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _057_ (
    .I0(p03[25]),
    .I1(p10[25]),
    .I2(p21[25]),
    .I3(p32[25]),
    .I4(key[89]),
    .O(z1[25])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _058_ (
    .I0(p03[26]),
    .I1(p10[26]),
    .I2(p21[26]),
    .I3(p32[26]),
    .I4(key[90]),
    .O(z1[26])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _059_ (
    .I0(p03[27]),
    .I1(p10[27]),
    .I2(p21[27]),
    .I3(p32[27]),
    .I4(key[91]),
    .O(z1[27])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _060_ (
    .I0(p03[28]),
    .I1(p10[28]),
    .I2(p21[28]),
    .I3(p32[28]),
    .I4(key[92]),
    .O(z1[28])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _061_ (
    .I0(p03[29]),
    .I1(p10[29]),
    .I2(p21[29]),
    .I3(p32[29]),
    .I4(key[93]),
    .O(z1[29])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _062_ (
    .I0(p03[30]),
    .I1(p10[30]),
    .I2(p21[30]),
    .I3(p32[30]),
    .I4(key[94]),
    .O(z1[30])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _063_ (
    .I0(p03[31]),
    .I1(p10[31]),
    .I2(p21[31]),
    .I3(p32[31]),
    .I4(key[95]),
    .O(z1[31])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _064_ (
    .I0(p02[0]),
    .I1(p13[0]),
    .I2(p20[0]),
    .I3(p31[0]),
    .I4(key[32]),
    .O(z2[0])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _065_ (
    .I0(p02[1]),
    .I1(p13[1]),
    .I2(p20[1]),
    .I3(p31[1]),
    .I4(key[33]),
    .O(z2[1])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _066_ (
    .I0(p02[2]),
    .I1(p13[2]),
    .I2(p20[2]),
    .I3(p31[2]),
    .I4(key[34]),
    .O(z2[2])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _067_ (
    .I0(p02[3]),
    .I1(p13[3]),
    .I2(p20[3]),
    .I3(p31[3]),
    .I4(key[35]),
    .O(z2[3])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _068_ (
    .I0(p02[4]),
    .I1(p13[4]),
    .I2(p20[4]),
    .I3(p31[4]),
    .I4(key[36]),
    .O(z2[4])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _069_ (
    .I0(p02[5]),
    .I1(p13[5]),
    .I2(p20[5]),
    .I3(p31[5]),
    .I4(key[37]),
    .O(z2[5])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _070_ (
    .I0(p02[6]),
    .I1(p13[6]),
    .I2(p20[6]),
    .I3(p31[6]),
    .I4(key[38]),
    .O(z2[6])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _071_ (
    .I0(p02[7]),
    .I1(p13[7]),
    .I2(p20[7]),
    .I3(p31[7]),
    .I4(key[39]),
    .O(z2[7])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _072_ (
    .I0(p02[8]),
    .I1(p13[8]),
    .I2(p20[8]),
    .I3(p31[8]),
    .I4(key[40]),
    .O(z2[8])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _073_ (
    .I0(p02[9]),
    .I1(p13[9]),
    .I2(p20[9]),
    .I3(p31[9]),
    .I4(key[41]),
    .O(z2[9])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _074_ (
    .I0(p02[10]),
    .I1(p13[10]),
    .I2(p20[10]),
    .I3(p31[10]),
    .I4(key[42]),
    .O(z2[10])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _075_ (
    .I0(p02[11]),
    .I1(p13[11]),
    .I2(p20[11]),
    .I3(p31[11]),
    .I4(key[43]),
    .O(z2[11])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _076_ (
    .I0(p02[12]),
    .I1(p13[12]),
    .I2(p20[12]),
    .I3(p31[12]),
    .I4(key[44]),
    .O(z2[12])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _077_ (
    .I0(p02[13]),
    .I1(p13[13]),
    .I2(p20[13]),
    .I3(p31[13]),
    .I4(key[45]),
    .O(z2[13])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _078_ (
    .I0(p02[14]),
    .I1(p13[14]),
    .I2(p20[14]),
    .I3(p31[14]),
    .I4(key[46]),
    .O(z2[14])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _079_ (
    .I0(p02[15]),
    .I1(p13[15]),
    .I2(p20[15]),
    .I3(p31[15]),
    .I4(key[47]),
    .O(z2[15])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _080_ (
    .I0(p02[16]),
    .I1(p13[16]),
    .I2(p20[16]),
    .I3(p31[16]),
    .I4(key[48]),
    .O(z2[16])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _081_ (
    .I0(p02[17]),
    .I1(p13[17]),
    .I2(p20[17]),
    .I3(p31[17]),
    .I4(key[49]),
    .O(z2[17])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _082_ (
    .I0(p02[18]),
    .I1(p13[18]),
    .I2(p20[18]),
    .I3(p31[18]),
    .I4(key[50]),
    .O(z2[18])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _083_ (
    .I0(p02[19]),
    .I1(p13[19]),
    .I2(p20[19]),
    .I3(p31[19]),
    .I4(key[51]),
    .O(z2[19])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _084_ (
    .I0(p02[20]),
    .I1(p13[20]),
    .I2(p20[20]),
    .I3(p31[20]),
    .I4(key[52]),
    .O(z2[20])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _085_ (
    .I0(p02[21]),
    .I1(p13[21]),
    .I2(p20[21]),
    .I3(p31[21]),
    .I4(key[53]),
    .O(z2[21])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _086_ (
    .I0(p02[22]),
    .I1(p13[22]),
    .I2(p20[22]),
    .I3(p31[22]),
    .I4(key[54]),
    .O(z2[22])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _087_ (
    .I0(p02[23]),
    .I1(p13[23]),
    .I2(p20[23]),
    .I3(p31[23]),
    .I4(key[55]),
    .O(z2[23])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _088_ (
    .I0(p02[24]),
    .I1(p13[24]),
    .I2(p20[24]),
    .I3(p31[24]),
    .I4(key[56]),
    .O(z2[24])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _089_ (
    .I0(p02[25]),
    .I1(p13[25]),
    .I2(p20[25]),
    .I3(p31[25]),
    .I4(key[57]),
    .O(z2[25])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _090_ (
    .I0(p02[26]),
    .I1(p13[26]),
    .I2(p20[26]),
    .I3(p31[26]),
    .I4(key[58]),
    .O(z2[26])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _091_ (
    .I0(p02[27]),
    .I1(p13[27]),
    .I2(p20[27]),
    .I3(p31[27]),
    .I4(key[59]),
    .O(z2[27])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _092_ (
    .I0(p02[28]),
    .I1(p13[28]),
    .I2(p20[28]),
    .I3(p31[28]),
    .I4(key[60]),
    .O(z2[28])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _093_ (
    .I0(p02[29]),
    .I1(p13[29]),
    .I2(p20[29]),
    .I3(p31[29]),
    .I4(key[61]),
    .O(z2[29])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _094_ (
    .I0(p02[30]),
    .I1(p13[30]),
    .I2(p20[30]),
    .I3(p31[30]),
    .I4(key[62]),
    .O(z2[30])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _095_ (
    .I0(p02[31]),
    .I1(p13[31]),
    .I2(p20[31]),
    .I3(p31[31]),
    .I4(key[63]),
    .O(z2[31])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _096_ (
    .I0(p01[0]),
    .I1(p12[0]),
    .I2(p23[0]),
    .I3(p30[0]),
    .I4(key[0]),
    .O(z3[0])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _097_ (
    .I0(p01[1]),
    .I1(p12[1]),
    .I2(p23[1]),
    .I3(p30[1]),
    .I4(key[1]),
    .O(z3[1])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _098_ (
    .I0(p01[2]),
    .I1(p12[2]),
    .I2(p23[2]),
    .I3(p30[2]),
    .I4(key[2]),
    .O(z3[2])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _099_ (
    .I0(p01[3]),
    .I1(p12[3]),
    .I2(p23[3]),
    .I3(p30[3]),
    .I4(key[3]),
    .O(z3[3])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _100_ (
    .I0(p01[4]),
    .I1(p12[4]),
    .I2(p23[4]),
    .I3(p30[4]),
    .I4(key[4]),
    .O(z3[4])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _101_ (
    .I0(p01[5]),
    .I1(p12[5]),
    .I2(p23[5]),
    .I3(p30[5]),
    .I4(key[5]),
    .O(z3[5])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _102_ (
    .I0(p01[6]),
    .I1(p12[6]),
    .I2(p23[6]),
    .I3(p30[6]),
    .I4(key[6]),
    .O(z3[6])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _103_ (
    .I0(p01[7]),
    .I1(p12[7]),
    .I2(p23[7]),
    .I3(p30[7]),
    .I4(key[7]),
    .O(z3[7])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _104_ (
    .I0(p01[8]),
    .I1(p12[8]),
    .I2(p23[8]),
    .I3(p30[8]),
    .I4(key[8]),
    .O(z3[8])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _105_ (
    .I0(p01[9]),
    .I1(p12[9]),
    .I2(p23[9]),
    .I3(p30[9]),
    .I4(key[9]),
    .O(z3[9])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _106_ (
    .I0(p01[10]),
    .I1(p12[10]),
    .I2(p23[10]),
    .I3(p30[10]),
    .I4(key[10]),
    .O(z3[10])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _107_ (
    .I0(p01[11]),
    .I1(p12[11]),
    .I2(p23[11]),
    .I3(p30[11]),
    .I4(key[11]),
    .O(z3[11])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _108_ (
    .I0(p01[12]),
    .I1(p12[12]),
    .I2(p23[12]),
    .I3(p30[12]),
    .I4(key[12]),
    .O(z3[12])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _109_ (
    .I0(p01[13]),
    .I1(p12[13]),
    .I2(p23[13]),
    .I3(p30[13]),
    .I4(key[13]),
    .O(z3[13])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _110_ (
    .I0(p01[14]),
    .I1(p12[14]),
    .I2(p23[14]),
    .I3(p30[14]),
    .I4(key[14]),
    .O(z3[14])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _111_ (
    .I0(p01[15]),
    .I1(p12[15]),
    .I2(p23[15]),
    .I3(p30[15]),
    .I4(key[15]),
    .O(z3[15])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _112_ (
    .I0(p01[16]),
    .I1(p12[16]),
    .I2(p23[16]),
    .I3(p30[16]),
    .I4(key[16]),
    .O(z3[16])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _113_ (
    .I0(p01[17]),
    .I1(p12[17]),
    .I2(p23[17]),
    .I3(p30[17]),
    .I4(key[17]),
    .O(z3[17])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _114_ (
    .I0(p01[18]),
    .I1(p12[18]),
    .I2(p23[18]),
    .I3(p30[18]),
    .I4(key[18]),
    .O(z3[18])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _115_ (
    .I0(p01[19]),
    .I1(p12[19]),
    .I2(p23[19]),
    .I3(p30[19]),
    .I4(key[19]),
    .O(z3[19])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _116_ (
    .I0(p01[20]),
    .I1(p12[20]),
    .I2(p23[20]),
    .I3(p30[20]),
    .I4(key[20]),
    .O(z3[20])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _117_ (
    .I0(p01[21]),
    .I1(p12[21]),
    .I2(p23[21]),
    .I3(p30[21]),
    .I4(key[21]),
    .O(z3[21])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _118_ (
    .I0(p01[22]),
    .I1(p12[22]),
    .I2(p23[22]),
    .I3(p30[22]),
    .I4(key[22]),
    .O(z3[22])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _119_ (
    .I0(p01[23]),
    .I1(p12[23]),
    .I2(p23[23]),
    .I3(p30[23]),
    .I4(key[23]),
    .O(z3[23])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _120_ (
    .I0(p01[24]),
    .I1(p12[24]),
    .I2(p23[24]),
    .I3(p30[24]),
    .I4(key[24]),
    .O(z3[24])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _121_ (
    .I0(p01[25]),
    .I1(p12[25]),
    .I2(p23[25]),
    .I3(p30[25]),
    .I4(key[25]),
    .O(z3[25])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _122_ (
    .I0(p01[26]),
    .I1(p12[26]),
    .I2(p23[26]),
    .I3(p30[26]),
    .I4(key[26]),
    .O(z3[26])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _123_ (
    .I0(p01[27]),
    .I1(p12[27]),
    .I2(p23[27]),
    .I3(p30[27]),
    .I4(key[27]),
    .O(z3[27])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _124_ (
    .I0(p01[28]),
    .I1(p12[28]),
    .I2(p23[28]),
    .I3(p30[28]),
    .I4(key[28]),
    .O(z3[28])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _125_ (
    .I0(p01[29]),
    .I1(p12[29]),
    .I2(p23[29]),
    .I3(p30[29]),
    .I4(key[29]),
    .O(z3[29])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _126_ (
    .I0(p01[30]),
    .I1(p12[30]),
    .I2(p23[30]),
    .I3(p30[30]),
    .I4(key[30]),
    .O(z3[30])
  );
LUT5  #(
    .INIT(32'd2523490710)
  ) _127_ (
    .I0(p01[31]),
    .I1(p12[31]),
    .I2(p23[31]),
    .I3(p30[31]),
    .I4(key[31]),
    .O(z3[31])
  );
FDRE  #(
    .INIT(1'hx)
  ) _128_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[0]),
    .Q(state_out[0]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _129_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[1]),
    .Q(state_out[1]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _130_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[2]),
    .Q(state_out[2]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _131_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[3]),
    .Q(state_out[3]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _132_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[4]),
    .Q(state_out[4]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _133_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[5]),
    .Q(state_out[5]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _134_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[6]),
    .Q(state_out[6]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _135_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[7]),
    .Q(state_out[7]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _136_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[8]),
    .Q(state_out[8]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _137_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[9]),
    .Q(state_out[9]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _138_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[10]),
    .Q(state_out[10]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _139_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[11]),
    .Q(state_out[11]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _140_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[12]),
    .Q(state_out[12]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _141_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[13]),
    .Q(state_out[13]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _142_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[14]),
    .Q(state_out[14]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _143_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[15]),
    .Q(state_out[15]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _144_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[16]),
    .Q(state_out[16]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _145_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[17]),
    .Q(state_out[17]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _146_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[18]),
    .Q(state_out[18]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _147_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[19]),
    .Q(state_out[19]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _148_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[20]),
    .Q(state_out[20]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _149_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[21]),
    .Q(state_out[21]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _150_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[22]),
    .Q(state_out[22]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _151_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[23]),
    .Q(state_out[23]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _152_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[24]),
    .Q(state_out[24]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _153_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[25]),
    .Q(state_out[25]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _154_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[26]),
    .Q(state_out[26]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _155_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[27]),
    .Q(state_out[27]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _156_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[28]),
    .Q(state_out[28]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _157_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[29]),
    .Q(state_out[29]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _158_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[30]),
    .Q(state_out[30]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _159_ (
    .C(clk),
    .CE(1'h1),
    .D(z3[31]),
    .Q(state_out[31]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _160_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[0]),
    .Q(state_out[32]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _161_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[1]),
    .Q(state_out[33]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _162_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[2]),
    .Q(state_out[34]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _163_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[3]),
    .Q(state_out[35]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _164_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[4]),
    .Q(state_out[36]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _165_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[5]),
    .Q(state_out[37]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _166_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[6]),
    .Q(state_out[38]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _167_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[7]),
    .Q(state_out[39]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _168_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[8]),
    .Q(state_out[40]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _169_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[9]),
    .Q(state_out[41]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _170_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[10]),
    .Q(state_out[42]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _171_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[11]),
    .Q(state_out[43]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _172_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[12]),
    .Q(state_out[44]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _173_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[13]),
    .Q(state_out[45]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _174_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[14]),
    .Q(state_out[46]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _175_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[15]),
    .Q(state_out[47]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _176_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[16]),
    .Q(state_out[48]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _177_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[17]),
    .Q(state_out[49]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _178_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[18]),
    .Q(state_out[50]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _179_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[19]),
    .Q(state_out[51]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _180_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[20]),
    .Q(state_out[52]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _181_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[21]),
    .Q(state_out[53]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _182_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[22]),
    .Q(state_out[54]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _183_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[23]),
    .Q(state_out[55]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _184_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[24]),
    .Q(state_out[56]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _185_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[25]),
    .Q(state_out[57]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _186_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[26]),
    .Q(state_out[58]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _187_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[27]),
    .Q(state_out[59]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _188_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[28]),
    .Q(state_out[60]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _189_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[29]),
    .Q(state_out[61]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _190_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[30]),
    .Q(state_out[62]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _191_ (
    .C(clk),
    .CE(1'h1),
    .D(z2[31]),
    .Q(state_out[63]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _192_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[0]),
    .Q(state_out[64]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _193_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[1]),
    .Q(state_out[65]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _194_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[2]),
    .Q(state_out[66]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _195_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[3]),
    .Q(state_out[67]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _196_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[4]),
    .Q(state_out[68]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _197_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[5]),
    .Q(state_out[69]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _198_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[6]),
    .Q(state_out[70]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _199_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[7]),
    .Q(state_out[71]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _200_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[8]),
    .Q(state_out[72]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _201_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[9]),
    .Q(state_out[73]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _202_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[10]),
    .Q(state_out[74]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _203_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[11]),
    .Q(state_out[75]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _204_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[12]),
    .Q(state_out[76]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _205_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[13]),
    .Q(state_out[77]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _206_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[14]),
    .Q(state_out[78]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _207_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[15]),
    .Q(state_out[79]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _208_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[16]),
    .Q(state_out[80]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _209_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[17]),
    .Q(state_out[81]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _210_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[18]),
    .Q(state_out[82]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _211_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[19]),
    .Q(state_out[83]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _212_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[20]),
    .Q(state_out[84]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _213_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[21]),
    .Q(state_out[85]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _214_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[22]),
    .Q(state_out[86]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _215_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[23]),
    .Q(state_out[87]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _216_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[24]),
    .Q(state_out[88]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _217_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[25]),
    .Q(state_out[89]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _218_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[26]),
    .Q(state_out[90]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _219_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[27]),
    .Q(state_out[91]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _220_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[28]),
    .Q(state_out[92]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _221_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[29]),
    .Q(state_out[93]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _222_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[30]),
    .Q(state_out[94]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _223_ (
    .C(clk),
    .CE(1'h1),
    .D(z1[31]),
    .Q(state_out[95]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _224_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[0]),
    .Q(state_out[96]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _225_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[1]),
    .Q(state_out[97]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _226_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[2]),
    .Q(state_out[98]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _227_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[3]),
    .Q(state_out[99]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _228_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[4]),
    .Q(state_out[100]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _229_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[5]),
    .Q(state_out[101]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _230_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[6]),
    .Q(state_out[102]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _231_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[7]),
    .Q(state_out[103]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _232_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[8]),
    .Q(state_out[104]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _233_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[9]),
    .Q(state_out[105]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _234_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[10]),
    .Q(state_out[106]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _235_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[11]),
    .Q(state_out[107]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _236_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[12]),
    .Q(state_out[108]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _237_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[13]),
    .Q(state_out[109]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _238_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[14]),
    .Q(state_out[110]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _239_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[15]),
    .Q(state_out[111]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _240_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[16]),
    .Q(state_out[112]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _241_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[17]),
    .Q(state_out[113]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _242_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[18]),
    .Q(state_out[114]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _243_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[19]),
    .Q(state_out[115]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _244_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[20]),
    .Q(state_out[116]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _245_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[21]),
    .Q(state_out[117]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _246_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[22]),
    .Q(state_out[118]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _247_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[23]),
    .Q(state_out[119]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _248_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[24]),
    .Q(state_out[120]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _249_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[25]),
    .Q(state_out[121]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _250_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[26]),
    .Q(state_out[122]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _251_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[27]),
    .Q(state_out[123]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _252_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[28]),
    .Q(state_out[124]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _253_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[29]),
    .Q(state_out[125]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _254_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[30]),
    .Q(state_out[126]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _255_ (
    .C(clk),
    .CE(1'h1),
    .D(z0[31]),
    .Q(state_out[127]),
    .R(1'h0)
  );
table_lookup  t0 (
    .clk(clk),
    .p0(p00),
    .p1(p01),
    .p2(p02),
    .p3(p03),
    .state(state_in[127:96])
  );
table_lookup  t1 (
    .clk(clk),
    .p0(p10),
    .p1(p11),
    .p2(p12),
    .p3(p13),
    .state(state_in[95:64])
  );
table_lookup  t2 (
    .clk(clk),
    .p0(p20),
    .p1(p21),
    .p2(p22),
    .p3(p23),
    .state(state_in[63:32])
  );
table_lookup  t3 (
    .clk(clk),
    .p0(p30),
    .p1(p31),
    .p2(p32),
    .p3(p33),
    .state(state_in[31:0])
  );
assign  k0 = key[127:96];
assign  k1 = key[95:64];
assign  k2 = key[63:32];
assign  k3 = key[31:0];
assign  s0 = state_in[127:96];
assign  s1 = state_in[95:64];
assign  s2 = state_in[63:32];
assign  s3 = state_in[31:0];
endmodule
