module S(clk,  in, out);
wire  _000_;
wire  _001_;
wire  _002_;
wire  _003_;
wire  _004_;
wire  _005_;
wire  _006_;
wire  _007_;
wire  _008_;
wire  _009_;
wire  _010_;
wire  _011_;
wire  _012_;
wire  _013_;
wire  _014_;
wire  _015_;
wire  _016_;
wire  _017_;
wire  _018_;
wire  _019_;
wire  _020_;
wire  _021_;
wire  _022_;
wire  _023_;
wire  _024_;
wire  _025_;
wire  _026_;
wire  _027_;
wire  _028_;
wire  _029_;
wire  _030_;
wire  _031_;
wire  _032_;
wire  _033_;
wire  _034_;
wire  _035_;
wire  _036_;
wire  _037_;
wire  _038_;
wire  _039_;
wire  _040_;
wire  _041_;
wire  _042_;
wire  _043_;
wire  _044_;
wire  _045_;
wire  _046_;
wire  _047_;
wire  [7:0] _048_;
input  clk;
input  [7:0] in;
output  [7:0] out;
LUT6  #(
    .INIT(64'h899a8190d169dd27)
  ) _049_ (
    .I0(in[6]),
    .I1(in[7]),
    .I2(in[4]),
    .I3(in[1]),
    .I4(in[5]),
    .I5(in[3]),
    .O(_002_)
  );
LUT6  #(
    .INIT(64'ha355cf0a13ce3106)
  ) _050_ (
    .I0(in[6]),
    .I1(in[7]),
    .I2(in[4]),
    .I3(in[1]),
    .I4(in[5]),
    .I5(in[3]),
    .O(_003_)
  );
MUXF7  _051_ (
    .I0(_002_),
    .I1(_003_),
    .O(_000_),
    .S(in[2])
  );
LUT6  #(
    .INIT(64'hab87bfaffab33162)
  ) _052_ (
    .I0(in[6]),
    .I1(in[7]),
    .I2(in[4]),
    .I3(in[1]),
    .I4(in[5]),
    .I5(in[3]),
    .O(_004_)
  );
LUT6  #(
    .INIT(64'h1d3c648f626b2595)
  ) _053_ (
    .I0(in[6]),
    .I1(in[7]),
    .I2(in[4]),
    .I3(in[1]),
    .I4(in[5]),
    .I5(in[3]),
    .O(_005_)
  );
MUXF7  _054_ (
    .I0(_004_),
    .I1(_005_),
    .O(_001_),
    .S(in[2])
  );
MUXF8  _055_ (
    .I0(_000_),
    .I1(_001_),
    .O(_048_[0]),
    .S(in[0])
  );
LUT6  #(
    .INIT(64'h710eb52f16199843)
  ) _056_ (
    .I0(in[5]),
    .I1(in[7]),
    .I2(in[6]),
    .I3(in[3]),
    .I4(in[4]),
    .I5(in[1]),
    .O(_008_)
  );
LUT6  #(
    .INIT(64'hafc971b356a5c137)
  ) _057_ (
    .I0(in[5]),
    .I1(in[7]),
    .I2(in[6]),
    .I3(in[3]),
    .I4(in[4]),
    .I5(in[1]),
    .O(_009_)
  );
MUXF7  _058_ (
    .I0(_008_),
    .I1(_009_),
    .O(_006_),
    .S(in[2])
  );
LUT6  #(
    .INIT(64'h8b62797b3e639c38)
  ) _059_ (
    .I0(in[5]),
    .I1(in[7]),
    .I2(in[6]),
    .I3(in[3]),
    .I4(in[4]),
    .I5(in[1]),
    .O(_010_)
  );
LUT6  #(
    .INIT(64'hf452c5442ec6115f)
  ) _060_ (
    .I0(in[5]),
    .I1(in[7]),
    .I2(in[6]),
    .I3(in[3]),
    .I4(in[4]),
    .I5(in[1]),
    .O(_011_)
  );
MUXF7  _061_ (
    .I0(_010_),
    .I1(_011_),
    .O(_007_),
    .S(in[2])
  );
MUXF8  _062_ (
    .I0(_006_),
    .I1(_007_),
    .O(_048_[1]),
    .S(in[0])
  );
LUT6  #(
    .INIT(64'h3d87b3b0530b8032)
  ) _063_ (
    .I0(in[0]),
    .I1(in[6]),
    .I2(in[7]),
    .I3(in[4]),
    .I4(in[5]),
    .I5(in[3]),
    .O(_014_)
  );
LUT6  #(
    .INIT(64'h9ae87bb3fa2b08f8)
  ) _064_ (
    .I0(in[0]),
    .I1(in[6]),
    .I2(in[7]),
    .I3(in[4]),
    .I4(in[5]),
    .I5(in[3]),
    .O(_015_)
  );
MUXF7  _065_ (
    .I0(_014_),
    .I1(_015_),
    .O(_012_),
    .S(in[2])
  );
LUT6  #(
    .INIT(64'hd05966f5b802fae5)
  ) _066_ (
    .I0(in[0]),
    .I1(in[6]),
    .I2(in[7]),
    .I3(in[4]),
    .I4(in[5]),
    .I5(in[3]),
    .O(_016_)
  );
LUT6  #(
    .INIT(64'h9296c80e19fbc1f3)
  ) _067_ (
    .I0(in[0]),
    .I1(in[6]),
    .I2(in[7]),
    .I3(in[4]),
    .I4(in[5]),
    .I5(in[3]),
    .O(_017_)
  );
MUXF7  _068_ (
    .I0(_016_),
    .I1(_017_),
    .O(_013_),
    .S(in[2])
  );
MUXF8  _069_ (
    .I0(_012_),
    .I1(_013_),
    .O(_048_[2]),
    .S(in[1])
  );
LUT6  #(
    .INIT(64'hc68322e46581880e)
  ) _070_ (
    .I0(in[7]),
    .I1(in[6]),
    .I2(in[5]),
    .I3(in[3]),
    .I4(in[4]),
    .I5(in[1]),
    .O(_020_)
  );
LUT6  #(
    .INIT(64'hade7cb6f8628ccdb)
  ) _071_ (
    .I0(in[7]),
    .I1(in[6]),
    .I2(in[5]),
    .I3(in[3]),
    .I4(in[4]),
    .I5(in[1]),
    .O(_021_)
  );
MUXF7  _072_ (
    .I0(_020_),
    .I1(_021_),
    .O(_018_),
    .S(in[0])
  );
LUT6  #(
    .INIT(64'hae60cf8517b98dae)
  ) _073_ (
    .I0(in[7]),
    .I1(in[6]),
    .I2(in[5]),
    .I3(in[3]),
    .I4(in[4]),
    .I5(in[1]),
    .O(_022_)
  );
LUT6  #(
    .INIT(64'h2ebee83066475ad5)
  ) _074_ (
    .I0(in[7]),
    .I1(in[6]),
    .I2(in[5]),
    .I3(in[3]),
    .I4(in[4]),
    .I5(in[1]),
    .O(_023_)
  );
MUXF7  _075_ (
    .I0(_022_),
    .I1(_023_),
    .O(_019_),
    .S(in[0])
  );
MUXF8  _076_ (
    .I0(_018_),
    .I1(_019_),
    .O(_048_[3]),
    .S(in[2])
  );
LUT6  #(
    .INIT(64'hf90a202aead99338)
  ) _077_ (
    .I0(in[6]),
    .I1(in[7]),
    .I2(in[5]),
    .I3(in[3]),
    .I4(in[0]),
    .I5(in[4]),
    .O(_026_)
  );
LUT6  #(
    .INIT(64'he473a5b1fd94711f)
  ) _078_ (
    .I0(in[6]),
    .I1(in[7]),
    .I2(in[5]),
    .I3(in[3]),
    .I4(in[0]),
    .I5(in[4]),
    .O(_027_)
  );
MUXF7  _079_ (
    .I0(_026_),
    .I1(_027_),
    .O(_024_),
    .S(in[2])
  );
LUT6  #(
    .INIT(64'h0e056e483ea30ed5)
  ) _080_ (
    .I0(in[6]),
    .I1(in[7]),
    .I2(in[5]),
    .I3(in[3]),
    .I4(in[0]),
    .I5(in[4]),
    .O(_028_)
  );
LUT6  #(
    .INIT(64'hbc33bb2ed5c4343a)
  ) _081_ (
    .I0(in[6]),
    .I1(in[7]),
    .I2(in[5]),
    .I3(in[3]),
    .I4(in[0]),
    .I5(in[4]),
    .O(_029_)
  );
MUXF7  _082_ (
    .I0(_028_),
    .I1(_029_),
    .O(_025_),
    .S(in[2])
  );
MUXF8  _083_ (
    .I0(_024_),
    .I1(_025_),
    .O(_048_[4]),
    .S(in[1])
  );
LUT6  #(
    .INIT(64'h9b792f252c2a79ad)
  ) _084_ (
    .I0(in[7]),
    .I1(in[5]),
    .I2(in[6]),
    .I3(in[1]),
    .I4(in[4]),
    .I5(in[3]),
    .O(_032_)
  );
LUT6  #(
    .INIT(64'h7d62df5639e067ed)
  ) _085_ (
    .I0(in[7]),
    .I1(in[5]),
    .I2(in[6]),
    .I3(in[1]),
    .I4(in[4]),
    .I5(in[3]),
    .O(_033_)
  );
MUXF7  _086_ (
    .I0(_032_),
    .I1(_033_),
    .O(_030_),
    .S(in[0])
  );
LUT6  #(
    .INIT(64'hcd8c9d1770936d85)
  ) _087_ (
    .I0(in[7]),
    .I1(in[5]),
    .I2(in[6]),
    .I3(in[1]),
    .I4(in[4]),
    .I5(in[3]),
    .O(_034_)
  );
LUT6  #(
    .INIT(64'h044d4b70c9921035)
  ) _088_ (
    .I0(in[7]),
    .I1(in[5]),
    .I2(in[6]),
    .I3(in[1]),
    .I4(in[4]),
    .I5(in[3]),
    .O(_035_)
  );
MUXF7  _089_ (
    .I0(_034_),
    .I1(_035_),
    .O(_031_),
    .S(in[0])
  );
MUXF8  _090_ (
    .I0(_030_),
    .I1(_031_),
    .O(_048_[5]),
    .S(in[2])
  );
LUT6  #(
    .INIT(64'hc4d0303d5fa6b827)
  ) _091_ (
    .I0(in[7]),
    .I1(in[0]),
    .I2(in[3]),
    .I3(in[6]),
    .I4(in[5]),
    .I5(in[1]),
    .O(_038_)
  );
LUT6  #(
    .INIT(64'h11ec2c0f21ae77e3)
  ) _092_ (
    .I0(in[7]),
    .I1(in[0]),
    .I2(in[3]),
    .I3(in[6]),
    .I4(in[5]),
    .I5(in[1]),
    .O(_039_)
  );
MUXF7  _093_ (
    .I0(_038_),
    .I1(_039_),
    .O(_036_),
    .S(in[4])
  );
LUT6  #(
    .INIT(64'h80ad09c7bf5264f7)
  ) _094_ (
    .I0(in[7]),
    .I1(in[0]),
    .I2(in[3]),
    .I3(in[6]),
    .I4(in[5]),
    .I5(in[1]),
    .O(_040_)
  );
LUT6  #(
    .INIT(64'h5e4256d5c8b8d6a5)
  ) _095_ (
    .I0(in[7]),
    .I1(in[0]),
    .I2(in[3]),
    .I3(in[6]),
    .I4(in[5]),
    .I5(in[1]),
    .O(_041_)
  );
MUXF7  _096_ (
    .I0(_040_),
    .I1(_041_),
    .O(_037_),
    .S(in[4])
  );
MUXF8  _097_ (
    .I0(_036_),
    .I1(_037_),
    .O(_048_[6]),
    .S(in[2])
  );
LUT6  #(
    .INIT(64'h994c6aea4c24de4e)
  ) _098_ (
    .I0(in[7]),
    .I1(in[5]),
    .I2(in[0]),
    .I3(in[6]),
    .I4(in[1]),
    .I5(in[3]),
    .O(_044_)
  );
LUT6  #(
    .INIT(64'h25dfd4315a61d8f9)
  ) _099_ (
    .I0(in[7]),
    .I1(in[5]),
    .I2(in[0]),
    .I3(in[6]),
    .I4(in[1]),
    .I5(in[3]),
    .O(_045_)
  );
MUXF7  _100_ (
    .I0(_044_),
    .I1(_045_),
    .O(_042_),
    .S(in[4])
  );
LUT6  #(
    .INIT(64'hf60938d9fa54a021)
  ) _101_ (
    .I0(in[7]),
    .I1(in[5]),
    .I2(in[0]),
    .I3(in[6]),
    .I4(in[1]),
    .I5(in[3]),
    .O(_046_)
  );
LUT6  #(
    .INIT(64'h7c3c6a1743f2dcc9)
  ) _102_ (
    .I0(in[7]),
    .I1(in[5]),
    .I2(in[0]),
    .I3(in[6]),
    .I4(in[1]),
    .I5(in[3]),
    .O(_047_)
  );
MUXF7  _103_ (
    .I0(_046_),
    .I1(_047_),
    .O(_043_),
    .S(in[4])
  );
MUXF8  _104_ (
    .I0(_042_),
    .I1(_043_),
    .O(_048_[7]),
    .S(in[2])
  );
FDRE  #(
    .INIT(1'hx)
  ) _105_ (
    .C(clk),
    .CE(1'h1),
    .D(_048_[0]),
    .Q(out[0]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _106_ (
    .C(clk),
    .CE(1'h1),
    .D(_048_[1]),
    .Q(out[1]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _107_ (
    .C(clk),
    .CE(1'h1),
    .D(_048_[2]),
    .Q(out[2]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _108_ (
    .C(clk),
    .CE(1'h1),
    .D(_048_[3]),
    .Q(out[3]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _109_ (
    .C(clk),
    .CE(1'h1),
    .D(_048_[4]),
    .Q(out[4]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _110_ (
    .C(clk),
    .CE(1'h1),
    .D(_048_[5]),
    .Q(out[5]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _111_ (
    .C(clk),
    .CE(1'h1),
    .D(_048_[6]),
    .Q(out[6]),
    .R(1'h0)
  );
FDRE  #(
    .INIT(1'hx)
  ) _112_ (
    .C(clk),
    .CE(1'h1),
    .D(_048_[7]),
    .Q(out[7]),
    .R(1'h0)
  );
endmodule
