module AES_Comp_InvMixColumns(x,  y);
wire  _000_;
wire  _001_;
wire  _002_;
wire  _003_;
wire  _004_;
wire  _005_;
wire  _006_;
wire  _007_;
wire  _008_;
wire  _009_;
wire  _010_;
wire  _011_;
wire  _012_;
wire  _013_;
wire  _014_;
wire  _015_;
wire  _016_;
wire  _017_;
wire  _018_;
wire  _019_;
wire  _020_;
wire  _021_;
wire  _022_;
wire  _023_;
wire  [1:0] _024_;
wire  [3:0] _025_;
wire  [4:0] _026_;
wire  [3:0] _027_;
wire  [5:0] _028_;
wire  [4:0] _029_;
wire  [2:0] _030_;
wire  [2:0] _031_;
wire  [4:0] _032_;
wire  [3:0] _033_;
wire  [5:0] _034_;
wire  [4:0] _035_;
wire  [2:0] _036_;
wire  [2:0] _037_;
wire  [2:0] _038_;
wire  [2:0] _039_;
wire  [7:0] a0;
wire  [7:0] a1;
wire  [7:0] a2;
wire  [7:0] a3;
input  [31:0] x;
wire  [31:0] x;
output  [31:0] y;
wire  [31:0] y;
LUT2  #(
    .INIT(4'h6)
  ) _040_ (
    .I0(_032_[0]),
    .I1(_033_[0]),
    .O(y[0])
  );
LUT5  #(
    .INIT(32'd1771476585)
  ) _041_ (
    .I0(x[24]),
    .I1(x[16]),
    .I2(x[31]),
    .I3(x[8]),
    .I4(x[7]),
    .O(_032_[0])
  );
LUT6  #(
    .INIT(64'h9669699669969669)
  ) _042_ (
    .I0(x[29]),
    .I1(x[21]),
    .I2(x[22]),
    .I3(x[13]),
    .I4(x[5]),
    .I5(x[6]),
    .O(_033_[0])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _043_ (
    .I0(_033_[0]),
    .I1(_033_[1]),
    .I2(_032_[1]),
    .I3(_032_[2]),
    .O(y[1])
  );
LUT6  #(
    .INIT(64'h9669699669969669)
  ) _044_ (
    .I0(x[24]),
    .I1(x[25]),
    .I2(x[17]),
    .I3(x[31]),
    .I4(x[9]),
    .I5(x[0]),
    .O(_000_)
  );
LUT6  #(
    .INIT(64'h6996966996696996)
  ) _045_ (
    .I0(x[24]),
    .I1(x[25]),
    .I2(x[17]),
    .I3(x[31]),
    .I4(x[9]),
    .I5(x[0]),
    .O(_001_)
  );
MUXF7  _046_ (
    .I0(_000_),
    .I1(_001_),
    .O(_033_[1]),
    .S(x[7])
  );
LUT5  #(
    .INIT(32'd1771476585)
  ) _047_ (
    .I0(x[22]),
    .I1(x[31]),
    .I2(x[14]),
    .I3(x[15]),
    .I4(x[7]),
    .O(_032_[1])
  );
LUT5  #(
    .INIT(32'd1771476585)
  ) _048_ (
    .I0(x[30]),
    .I1(x[31]),
    .I2(x[23]),
    .I3(x[15]),
    .I4(x[6]),
    .O(_032_[2])
  );
LUT5  #(
    .INIT(32'd1771476585)
  ) _049_ (
    .I0(_032_[0]),
    .I1(_032_[1]),
    .I2(_032_[2]),
    .I3(_032_[3]),
    .I4(_034_[3]),
    .O(y[2])
  );
LUT5  #(
    .INIT(32'd1771476585)
  ) _050_ (
    .I0(x[24]),
    .I1(x[23]),
    .I2(x[8]),
    .I3(x[15]),
    .I4(x[0]),
    .O(_032_[3])
  );
LUT5  #(
    .INIT(32'd1771476585)
  ) _051_ (
    .I0(x[25]),
    .I1(x[26]),
    .I2(x[18]),
    .I3(x[10]),
    .I4(x[1]),
    .O(_034_[3])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _052_ (
    .I0(_033_[0]),
    .I1(_033_[1]),
    .I2(_033_[2]),
    .I3(_035_[2]),
    .O(y[3])
  );
LUT6  #(
    .INIT(64'h9669699669969669)
  ) _053_ (
    .I0(x[16]),
    .I1(x[25]),
    .I2(x[23]),
    .I3(x[8]),
    .I4(x[9]),
    .I5(x[15]),
    .O(_002_)
  );
LUT6  #(
    .INIT(64'h6996966996696996)
  ) _054_ (
    .I0(x[16]),
    .I1(x[25]),
    .I2(x[23]),
    .I3(x[8]),
    .I4(x[9]),
    .I5(x[15]),
    .O(_003_)
  );
MUXF7  _055_ (
    .I0(_002_),
    .I1(_003_),
    .O(_033_[2]),
    .S(x[1])
  );
LUT6  #(
    .INIT(64'h9669699669969669)
  ) _056_ (
    .I0(x[26]),
    .I1(x[27]),
    .I2(x[19]),
    .I3(x[31]),
    .I4(x[11]),
    .I5(x[2]),
    .O(_004_)
  );
LUT6  #(
    .INIT(64'h6996966996696996)
  ) _057_ (
    .I0(x[26]),
    .I1(x[27]),
    .I2(x[19]),
    .I3(x[31]),
    .I4(x[11]),
    .I5(x[2]),
    .O(_005_)
  );
MUXF7  _058_ (
    .I0(_004_),
    .I1(_005_),
    .O(_035_[2]),
    .S(x[7])
  );
LUT6  #(
    .INIT(64'h6996966996696996)
  ) _059_ (
    .I0(_033_[0]),
    .I1(_032_[1]),
    .I2(_032_[2]),
    .I3(_034_[3]),
    .I4(_032_[4]),
    .I5(_036_[1]),
    .O(y[4])
  );
LUT5  #(
    .INIT(32'd1771476585)
  ) _060_ (
    .I0(x[17]),
    .I1(x[26]),
    .I2(x[9]),
    .I3(x[10]),
    .I4(x[2]),
    .O(_032_[4])
  );
LUT6  #(
    .INIT(64'h9669699669969669)
  ) _061_ (
    .I0(x[27]),
    .I1(x[28]),
    .I2(x[20]),
    .I3(x[31]),
    .I4(x[12]),
    .I5(x[3]),
    .O(_006_)
  );
LUT6  #(
    .INIT(64'h6996966996696996)
  ) _062_ (
    .I0(x[27]),
    .I1(x[28]),
    .I2(x[20]),
    .I3(x[31]),
    .I4(x[12]),
    .I5(x[3]),
    .O(_007_)
  );
MUXF7  _063_ (
    .I0(_006_),
    .I1(_007_),
    .O(_036_[1]),
    .S(x[7])
  );
LUT5  #(
    .INIT(32'd1771476585)
  ) _064_ (
    .I0(_032_[1]),
    .I1(_032_[2]),
    .I2(_035_[2]),
    .I3(_033_[3]),
    .I4(_037_[1]),
    .O(y[5])
  );
LUT6  #(
    .INIT(64'h9669699669969669)
  ) _065_ (
    .I0(x[18]),
    .I1(x[27]),
    .I2(x[23]),
    .I3(x[10]),
    .I4(x[11]),
    .I5(x[15]),
    .O(_008_)
  );
LUT6  #(
    .INIT(64'h6996966996696996)
  ) _066_ (
    .I0(x[18]),
    .I1(x[27]),
    .I2(x[23]),
    .I3(x[10]),
    .I4(x[11]),
    .I5(x[15]),
    .O(_009_)
  );
MUXF7  _067_ (
    .I0(_008_),
    .I1(_009_),
    .O(_033_[3]),
    .S(x[3])
  );
LUT5  #(
    .INIT(32'd1771476585)
  ) _068_ (
    .I0(x[28]),
    .I1(x[29]),
    .I2(x[21]),
    .I3(x[13]),
    .I4(x[4]),
    .O(_037_[1])
  );
LUT3  #(
    .INIT(8'h69)
  ) _069_ (
    .I0(_038_[0]),
    .I1(_036_[1]),
    .I2(_034_[5]),
    .O(y[6])
  );
LUT5  #(
    .INIT(32'd1771476585)
  ) _070_ (
    .I0(x[29]),
    .I1(x[30]),
    .I2(x[22]),
    .I3(x[14]),
    .I4(x[5]),
    .O(_038_[0])
  );
LUT6  #(
    .INIT(64'h9669699669969669)
  ) _071_ (
    .I0(x[19]),
    .I1(x[28]),
    .I2(x[23]),
    .I3(x[11]),
    .I4(x[12]),
    .I5(x[15]),
    .O(_010_)
  );
LUT6  #(
    .INIT(64'h6996966996696996)
  ) _072_ (
    .I0(x[19]),
    .I1(x[28]),
    .I2(x[23]),
    .I3(x[11]),
    .I4(x[12]),
    .I5(x[15]),
    .O(_011_)
  );
MUXF7  _073_ (
    .I0(_010_),
    .I1(_011_),
    .O(_034_[5]),
    .S(x[4])
  );
LUT3  #(
    .INIT(8'h69)
  ) _074_ (
    .I0(_032_[2]),
    .I1(_037_[1]),
    .I2(_035_[4]),
    .O(y[7])
  );
LUT5  #(
    .INIT(32'd1771476585)
  ) _075_ (
    .I0(x[20]),
    .I1(x[29]),
    .I2(x[12]),
    .I3(x[13]),
    .I4(x[5]),
    .O(_035_[4])
  );
LUT2  #(
    .INIT(4'h6)
  ) _076_ (
    .I0(_026_[0]),
    .I1(_024_[0]),
    .O(y[8])
  );
LUT5  #(
    .INIT(32'd1771476585)
  ) _077_ (
    .I0(x[24]),
    .I1(x[16]),
    .I2(x[15]),
    .I3(x[0]),
    .I4(x[7]),
    .O(_026_[0])
  );
LUT6  #(
    .INIT(64'h9669699669969669)
  ) _078_ (
    .I0(x[29]),
    .I1(x[21]),
    .I2(x[30]),
    .I3(x[13]),
    .I4(x[14]),
    .I5(x[5]),
    .O(_024_[0])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _079_ (
    .I0(_024_[0]),
    .I1(_027_[1]),
    .I2(_025_[1]),
    .I3(_025_[2]),
    .O(y[9])
  );
LUT6  #(
    .INIT(64'h9669699669969669)
  ) _080_ (
    .I0(x[25]),
    .I1(x[17]),
    .I2(x[8]),
    .I3(x[15]),
    .I4(x[0]),
    .I5(x[1]),
    .O(_012_)
  );
LUT6  #(
    .INIT(64'h6996966996696996)
  ) _081_ (
    .I0(x[25]),
    .I1(x[17]),
    .I2(x[8]),
    .I3(x[15]),
    .I4(x[0]),
    .I5(x[1]),
    .O(_013_)
  );
MUXF7  _082_ (
    .I0(_012_),
    .I1(_013_),
    .O(_027_[1]),
    .S(x[7])
  );
LUT5  #(
    .INIT(32'd1771476585)
  ) _083_ (
    .I0(x[30]),
    .I1(x[22]),
    .I2(x[23]),
    .I3(x[15]),
    .I4(x[7]),
    .O(_025_[1])
  );
LUT5  #(
    .INIT(32'd1771476585)
  ) _084_ (
    .I0(x[31]),
    .I1(x[23]),
    .I2(x[14]),
    .I3(x[6]),
    .I4(x[7]),
    .O(_025_[2])
  );
LUT5  #(
    .INIT(32'd1771476585)
  ) _085_ (
    .I0(_026_[0]),
    .I1(_025_[1]),
    .I2(_025_[2]),
    .I3(_024_[1]),
    .I4(_028_[3]),
    .O(y[10])
  );
LUT5  #(
    .INIT(32'd1771476585)
  ) _086_ (
    .I0(x[16]),
    .I1(x[31]),
    .I2(x[23]),
    .I3(x[8]),
    .I4(x[0]),
    .O(_024_[1])
  );
LUT5  #(
    .INIT(32'd1771476585)
  ) _087_ (
    .I0(x[26]),
    .I1(x[18]),
    .I2(x[9]),
    .I3(x[1]),
    .I4(x[2]),
    .O(_028_[3])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _088_ (
    .I0(_024_[0]),
    .I1(_027_[1]),
    .I2(_025_[3]),
    .I3(_029_[2]),
    .O(y[11])
  );
LUT6  #(
    .INIT(64'h9669699669969669)
  ) _089_ (
    .I0(x[24]),
    .I1(x[16]),
    .I2(x[17]),
    .I3(x[31]),
    .I4(x[23]),
    .I5(x[9]),
    .O(_014_)
  );
LUT6  #(
    .INIT(64'h6996966996696996)
  ) _090_ (
    .I0(x[24]),
    .I1(x[16]),
    .I2(x[17]),
    .I3(x[31]),
    .I4(x[23]),
    .I5(x[9]),
    .O(_015_)
  );
MUXF7  _091_ (
    .I0(_014_),
    .I1(_015_),
    .O(_025_[3]),
    .S(x[1])
  );
LUT6  #(
    .INIT(64'h9669699669969669)
  ) _092_ (
    .I0(x[27]),
    .I1(x[19]),
    .I2(x[10]),
    .I3(x[15]),
    .I4(x[2]),
    .I5(x[3]),
    .O(_016_)
  );
LUT6  #(
    .INIT(64'h6996966996696996)
  ) _093_ (
    .I0(x[27]),
    .I1(x[19]),
    .I2(x[10]),
    .I3(x[15]),
    .I4(x[2]),
    .I5(x[3]),
    .O(_017_)
  );
MUXF7  _094_ (
    .I0(_016_),
    .I1(_017_),
    .O(_029_[2]),
    .S(x[7])
  );
LUT6  #(
    .INIT(64'h6996966996696996)
  ) _095_ (
    .I0(_024_[0]),
    .I1(_025_[1]),
    .I2(_025_[2]),
    .I3(_028_[3]),
    .I4(_026_[4]),
    .I5(_030_[1]),
    .O(y[12])
  );
LUT5  #(
    .INIT(32'd1771476585)
  ) _096_ (
    .I0(x[25]),
    .I1(x[17]),
    .I2(x[18]),
    .I3(x[10]),
    .I4(x[2]),
    .O(_026_[4])
  );
LUT6  #(
    .INIT(64'h9669699669969669)
  ) _097_ (
    .I0(x[28]),
    .I1(x[20]),
    .I2(x[11]),
    .I3(x[15]),
    .I4(x[3]),
    .I5(x[4]),
    .O(_018_)
  );
LUT6  #(
    .INIT(64'h6996966996696996)
  ) _098_ (
    .I0(x[28]),
    .I1(x[20]),
    .I2(x[11]),
    .I3(x[15]),
    .I4(x[3]),
    .I5(x[4]),
    .O(_019_)
  );
MUXF7  _099_ (
    .I0(_018_),
    .I1(_019_),
    .O(_030_[1]),
    .S(x[7])
  );
LUT5  #(
    .INIT(32'd1771476585)
  ) _100_ (
    .I0(_025_[1]),
    .I1(_025_[2]),
    .I2(_029_[2]),
    .I3(_027_[3]),
    .I4(_031_[1]),
    .O(y[13])
  );
LUT6  #(
    .INIT(64'h9669699669969669)
  ) _101_ (
    .I0(x[26]),
    .I1(x[18]),
    .I2(x[19]),
    .I3(x[31]),
    .I4(x[23]),
    .I5(x[11]),
    .O(_020_)
  );
LUT6  #(
    .INIT(64'h6996966996696996)
  ) _102_ (
    .I0(x[26]),
    .I1(x[18]),
    .I2(x[19]),
    .I3(x[31]),
    .I4(x[23]),
    .I5(x[11]),
    .O(_021_)
  );
MUXF7  _103_ (
    .I0(_020_),
    .I1(_021_),
    .O(_027_[3]),
    .S(x[3])
  );
LUT5  #(
    .INIT(32'd1771476585)
  ) _104_ (
    .I0(x[29]),
    .I1(x[21]),
    .I2(x[12]),
    .I3(x[4]),
    .I4(x[5]),
    .O(_031_[1])
  );
LUT3  #(
    .INIT(8'h69)
  ) _105_ (
    .I0(_039_[0]),
    .I1(_030_[1]),
    .I2(_028_[5]),
    .O(y[14])
  );
LUT5  #(
    .INIT(32'd1771476585)
  ) _106_ (
    .I0(x[30]),
    .I1(x[22]),
    .I2(x[13]),
    .I3(x[5]),
    .I4(x[6]),
    .O(_039_[0])
  );
LUT6  #(
    .INIT(64'h9669699669969669)
  ) _107_ (
    .I0(x[27]),
    .I1(x[19]),
    .I2(x[20]),
    .I3(x[31]),
    .I4(x[23]),
    .I5(x[12]),
    .O(_022_)
  );
LUT6  #(
    .INIT(64'h6996966996696996)
  ) _108_ (
    .I0(x[27]),
    .I1(x[19]),
    .I2(x[20]),
    .I3(x[31]),
    .I4(x[23]),
    .I5(x[12]),
    .O(_023_)
  );
MUXF7  _109_ (
    .I0(_022_),
    .I1(_023_),
    .O(_028_[5]),
    .S(x[4])
  );
LUT3  #(
    .INIT(8'h69)
  ) _110_ (
    .I0(_025_[2]),
    .I1(_031_[1]),
    .I2(_029_[4]),
    .O(y[15])
  );
LUT5  #(
    .INIT(32'd1771476585)
  ) _111_ (
    .I0(x[28]),
    .I1(x[20]),
    .I2(x[21]),
    .I3(x[13]),
    .I4(x[5]),
    .O(_029_[4])
  );
LUT2  #(
    .INIT(4'h6)
  ) _112_ (
    .I0(_033_[0]),
    .I1(_032_[3]),
    .O(y[16])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _113_ (
    .I0(_033_[0]),
    .I1(_032_[1]),
    .I2(_032_[2]),
    .I3(_033_[2]),
    .O(y[17])
  );
LUT5  #(
    .INIT(32'd1771476585)
  ) _114_ (
    .I0(_032_[0]),
    .I1(_032_[1]),
    .I2(_032_[2]),
    .I3(_032_[3]),
    .I4(_032_[4]),
    .O(y[18])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _115_ (
    .I0(_033_[0]),
    .I1(_033_[1]),
    .I2(_033_[2]),
    .I3(_033_[3]),
    .O(y[19])
  );
LUT6  #(
    .INIT(64'h6996966996696996)
  ) _116_ (
    .I0(_033_[0]),
    .I1(_032_[1]),
    .I2(_032_[2]),
    .I3(_034_[3]),
    .I4(_032_[4]),
    .I5(_034_[5]),
    .O(y[20])
  );
LUT5  #(
    .INIT(32'd1771476585)
  ) _117_ (
    .I0(_032_[1]),
    .I1(_032_[2]),
    .I2(_035_[2]),
    .I3(_033_[3]),
    .I4(_035_[4]),
    .O(y[21])
  );
LUT3  #(
    .INIT(8'h69)
  ) _118_ (
    .I0(_036_[0]),
    .I1(_036_[1]),
    .I2(_034_[5]),
    .O(y[22])
  );
LUT5  #(
    .INIT(32'd1771476585)
  ) _119_ (
    .I0(x[21]),
    .I1(x[30]),
    .I2(x[13]),
    .I3(x[14]),
    .I4(x[6]),
    .O(_036_[0])
  );
LUT3  #(
    .INIT(8'h69)
  ) _120_ (
    .I0(_032_[1]),
    .I1(_037_[1]),
    .I2(_035_[4]),
    .O(y[23])
  );
LUT2  #(
    .INIT(4'h6)
  ) _121_ (
    .I0(_024_[0]),
    .I1(_024_[1]),
    .O(y[24])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _122_ (
    .I0(_024_[0]),
    .I1(_025_[1]),
    .I2(_025_[2]),
    .I3(_025_[3]),
    .O(y[25])
  );
LUT5  #(
    .INIT(32'd1771476585)
  ) _123_ (
    .I0(_026_[0]),
    .I1(_025_[1]),
    .I2(_025_[2]),
    .I3(_024_[1]),
    .I4(_026_[4]),
    .O(y[26])
  );
LUT4  #(
    .INIT(16'h6996)
  ) _124_ (
    .I0(_024_[0]),
    .I1(_027_[1]),
    .I2(_025_[3]),
    .I3(_027_[3]),
    .O(y[27])
  );
LUT6  #(
    .INIT(64'h6996966996696996)
  ) _125_ (
    .I0(_024_[0]),
    .I1(_025_[1]),
    .I2(_025_[2]),
    .I3(_028_[3]),
    .I4(_026_[4]),
    .I5(_028_[5]),
    .O(y[28])
  );
LUT5  #(
    .INIT(32'd1771476585)
  ) _126_ (
    .I0(_025_[1]),
    .I1(_025_[2]),
    .I2(_029_[2]),
    .I3(_027_[3]),
    .I4(_029_[4]),
    .O(y[29])
  );
LUT3  #(
    .INIT(8'h69)
  ) _127_ (
    .I0(_030_[0]),
    .I1(_030_[1]),
    .I2(_028_[5]),
    .O(y[30])
  );
LUT5  #(
    .INIT(32'd1771476585)
  ) _128_ (
    .I0(x[29]),
    .I1(x[21]),
    .I2(x[22]),
    .I3(x[14]),
    .I4(x[6]),
    .O(_030_[0])
  );
LUT3  #(
    .INIT(8'h69)
  ) _129_ (
    .I0(_025_[1]),
    .I1(_031_[1]),
    .I2(_029_[4]),
    .O(y[31])
  );
assign  { _034_[4], _034_[2:0] } = { _032_[4], _032_[2:1], _033_[0] };
assign  _036_[2] = _034_[5];
assign  { _028_[4], _028_[2:0] } = { _026_[4], _025_[2:1], _024_[0] };
assign  { _027_[2], _027_[0] } = { _025_[3], _024_[0] };
assign  _039_[2:1] = { _028_[5], _030_[1] };
assign  { _031_[2], _031_[0] } = { _029_[4], _025_[1] };
assign  { _037_[2], _037_[0] } = { _035_[4], _032_[1] };
assign  _026_[3:1] = { _024_[1], _025_[2:1] };
assign  { _035_[3], _035_[1:0] } = { _033_[3], _032_[2:1] };
assign  _030_[2] = _028_[5];
assign  _025_[0] = _024_[0];
assign  { _029_[3], _029_[1:0] } = { _027_[3], _025_[2:1] };
assign  _038_[2:1] = { _034_[5], _036_[1] };
assign  a0 = x[7:0];
assign  a1 = x[15:8];
assign  a2 = x[23:16];
assign  a3 = x[31:24];
endmodule
