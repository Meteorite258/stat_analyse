module AES_Comp_GFinvComp(x,  y);
wire  _000_;
wire  _001_;
wire  _002_;
wire  _003_;
wire  _004_;
wire  _005_;
wire  _006_;
wire  _007_;
wire  _008_;
wire  _009_;
wire  _010_;
wire  _011_;
wire  _012_;
wire  _013_;
wire  _014_;
wire  _015_;
wire  _016_;
wire  _017_;
wire  _018_;
wire  _019_;
wire  _020_;
wire  _021_;
wire  _022_;
wire  _023_;
wire  _024_;
wire  _025_;
wire  _026_;
wire  _027_;
wire  _028_;
wire  _029_;
wire  _030_;
wire  _031_;
wire  _032_;
wire  _033_;
wire  _034_;
wire  _035_;
wire  _036_;
wire  _037_;
wire  _038_;
wire  _039_;
wire  _040_;
wire  _041_;
wire  _042_;
wire  _043_;
wire  _044_;
wire  _045_;
wire  _046_;
wire  _047_;
wire  [8:0] da;
wire  [8:0] db;
input  [7:0] x;
wire  [7:0] x;
output  [7:0] y;
wire  [7:0] y;
LUT6  #(
    .INIT(64'hb5f6225d259e3d86)
  ) _048_ (
    .I0(x[0]),
    .I1(x[1]),
    .I2(x[3]),
    .I3(x[4]),
    .I4(x[6]),
    .I5(x[2]),
    .O(_002_)
  );
LUT6  #(
    .INIT(64'hd75b6c3f520074e9)
  ) _049_ (
    .I0(x[0]),
    .I1(x[1]),
    .I2(x[3]),
    .I3(x[4]),
    .I4(x[6]),
    .I5(x[2]),
    .O(_003_)
  );
MUXF7  _050_ (
    .I0(_002_),
    .I1(_003_),
    .O(_000_),
    .S(x[5])
  );
LUT6  #(
    .INIT(64'h984e5dd4737940eb)
  ) _051_ (
    .I0(x[0]),
    .I1(x[1]),
    .I2(x[3]),
    .I3(x[4]),
    .I4(x[6]),
    .I5(x[2]),
    .O(_004_)
  );
LUT6  #(
    .INIT(64'h433a42dab0c829b9)
  ) _052_ (
    .I0(x[0]),
    .I1(x[1]),
    .I2(x[3]),
    .I3(x[4]),
    .I4(x[6]),
    .I5(x[2]),
    .O(_005_)
  );
MUXF7  _053_ (
    .I0(_004_),
    .I1(_005_),
    .O(_001_),
    .S(x[5])
  );
MUXF8  _054_ (
    .I0(_000_),
    .I1(_001_),
    .O(y[0]),
    .S(x[7])
  );
LUT6  #(
    .INIT(64'hef53544bdac82b9c)
  ) _055_ (
    .I0(x[0]),
    .I1(x[1]),
    .I2(x[2]),
    .I3(x[3]),
    .I4(x[4]),
    .I5(x[5]),
    .O(_008_)
  );
LUT6  #(
    .INIT(64'ha652d2357580de83)
  ) _056_ (
    .I0(x[0]),
    .I1(x[1]),
    .I2(x[2]),
    .I3(x[3]),
    .I4(x[4]),
    .I5(x[5]),
    .O(_009_)
  );
MUXF7  _057_ (
    .I0(_008_),
    .I1(_009_),
    .O(_006_),
    .S(x[6])
  );
LUT6  #(
    .INIT(64'h079049799db43cfe)
  ) _058_ (
    .I0(x[0]),
    .I1(x[1]),
    .I2(x[2]),
    .I3(x[3]),
    .I4(x[4]),
    .I5(x[5]),
    .O(_010_)
  );
LUT6  #(
    .INIT(64'h76b38b904483e8b7)
  ) _059_ (
    .I0(x[0]),
    .I1(x[1]),
    .I2(x[2]),
    .I3(x[3]),
    .I4(x[4]),
    .I5(x[5]),
    .O(_011_)
  );
MUXF7  _060_ (
    .I0(_010_),
    .I1(_011_),
    .O(_007_),
    .S(x[6])
  );
MUXF8  _061_ (
    .I0(_006_),
    .I1(_007_),
    .O(y[1]),
    .S(x[7])
  );
LUT6  #(
    .INIT(64'hf47b3ad372fca544)
  ) _062_ (
    .I0(x[1]),
    .I1(x[2]),
    .I2(x[0]),
    .I3(x[4]),
    .I4(x[3]),
    .I5(x[6]),
    .O(_014_)
  );
LUT6  #(
    .INIT(64'h26bf6b23caab1879)
  ) _063_ (
    .I0(x[1]),
    .I1(x[2]),
    .I2(x[0]),
    .I3(x[4]),
    .I4(x[3]),
    .I5(x[6]),
    .O(_015_)
  );
MUXF7  _064_ (
    .I0(_014_),
    .I1(_015_),
    .O(_012_),
    .S(x[5])
  );
LUT6  #(
    .INIT(64'hbd03bc9de09250ce)
  ) _065_ (
    .I0(x[1]),
    .I1(x[2]),
    .I2(x[0]),
    .I3(x[4]),
    .I4(x[3]),
    .I5(x[6]),
    .O(_016_)
  );
LUT6  #(
    .INIT(64'h2983d21193f05b42)
  ) _066_ (
    .I0(x[1]),
    .I1(x[2]),
    .I2(x[0]),
    .I3(x[4]),
    .I4(x[3]),
    .I5(x[6]),
    .O(_017_)
  );
MUXF7  _067_ (
    .I0(_016_),
    .I1(_017_),
    .O(_013_),
    .S(x[5])
  );
MUXF8  _068_ (
    .I0(_012_),
    .I1(_013_),
    .O(y[2]),
    .S(x[7])
  );
LUT6  #(
    .INIT(64'hdac7e52588e263f0)
  ) _069_ (
    .I0(x[1]),
    .I1(x[0]),
    .I2(x[2]),
    .I3(x[3]),
    .I4(x[4]),
    .I5(x[5]),
    .O(_020_)
  );
LUT6  #(
    .INIT(64'h90437dd6568a9d03)
  ) _070_ (
    .I0(x[1]),
    .I1(x[0]),
    .I2(x[2]),
    .I3(x[3]),
    .I4(x[4]),
    .I5(x[5]),
    .O(_021_)
  );
MUXF7  _071_ (
    .I0(_020_),
    .I1(_021_),
    .O(_018_),
    .S(x[6])
  );
LUT6  #(
    .INIT(64'hf0dd687eca1df6ab)
  ) _072_ (
    .I0(x[1]),
    .I1(x[0]),
    .I2(x[2]),
    .I3(x[3]),
    .I4(x[4]),
    .I5(x[5]),
    .O(_022_)
  );
LUT6  #(
    .INIT(64'h62684262ba4baf48)
  ) _073_ (
    .I0(x[1]),
    .I1(x[0]),
    .I2(x[2]),
    .I3(x[3]),
    .I4(x[4]),
    .I5(x[5]),
    .O(_023_)
  );
MUXF7  _074_ (
    .I0(_022_),
    .I1(_023_),
    .O(_019_),
    .S(x[6])
  );
MUXF8  _075_ (
    .I0(_018_),
    .I1(_019_),
    .O(y[3]),
    .S(x[7])
  );
LUT6  #(
    .INIT(64'ha5ff303366880000)
  ) _076_ (
    .I0(x[0]),
    .I1(x[1]),
    .I2(x[2]),
    .I3(x[3]),
    .I4(x[6]),
    .I5(x[4]),
    .O(_026_)
  );
LUT6  #(
    .INIT(64'ha335b478d99d9595)
  ) _077_ (
    .I0(x[0]),
    .I1(x[1]),
    .I2(x[2]),
    .I3(x[3]),
    .I4(x[6]),
    .I5(x[4]),
    .O(_027_)
  );
MUXF7  _078_ (
    .I0(_026_),
    .I1(_027_),
    .O(_024_),
    .S(x[7])
  );
LUT6  #(
    .INIT(64'h7e3c09f655bef50f)
  ) _079_ (
    .I0(x[0]),
    .I1(x[1]),
    .I2(x[2]),
    .I3(x[3]),
    .I4(x[6]),
    .I5(x[4]),
    .O(_028_)
  );
LUT6  #(
    .INIT(64'h47e20b0d16947dd7)
  ) _080_ (
    .I0(x[0]),
    .I1(x[1]),
    .I2(x[2]),
    .I3(x[3]),
    .I4(x[6]),
    .I5(x[4]),
    .O(_029_)
  );
MUXF7  _081_ (
    .I0(_028_),
    .I1(_029_),
    .O(_025_),
    .S(x[7])
  );
MUXF8  _082_ (
    .I0(_024_),
    .I1(_025_),
    .O(y[4]),
    .S(x[5])
  );
LUT6  #(
    .INIT(64'h9f6f0555c2c20000)
  ) _083_ (
    .I0(x[0]),
    .I1(x[1]),
    .I2(x[2]),
    .I3(x[3]),
    .I4(x[7]),
    .I5(x[5]),
    .O(_032_)
  );
LUT6  #(
    .INIT(64'h979e90ffe5da3f0c)
  ) _084_ (
    .I0(x[0]),
    .I1(x[1]),
    .I2(x[2]),
    .I3(x[3]),
    .I4(x[7]),
    .I5(x[5]),
    .O(_033_)
  );
MUXF7  _085_ (
    .I0(_032_),
    .I1(_033_),
    .O(_030_),
    .S(x[4])
  );
LUT6  #(
    .INIT(64'h8d725569933933bb)
  ) _086_ (
    .I0(x[0]),
    .I1(x[1]),
    .I2(x[2]),
    .I3(x[3]),
    .I4(x[7]),
    .I5(x[5]),
    .O(_034_)
  );
LUT6  #(
    .INIT(64'hbbddc318700bde84)
  ) _087_ (
    .I0(x[0]),
    .I1(x[1]),
    .I2(x[2]),
    .I3(x[3]),
    .I4(x[7]),
    .I5(x[5]),
    .O(_035_)
  );
MUXF7  _088_ (
    .I0(_034_),
    .I1(_035_),
    .O(_031_),
    .S(x[4])
  );
MUXF8  _089_ (
    .I0(_030_),
    .I1(_031_),
    .O(y[5]),
    .S(x[6])
  );
LUT6  #(
    .INIT(64'h4d8e30fcf9f90000)
  ) _090_ (
    .I0(x[3]),
    .I1(x[0]),
    .I2(x[2]),
    .I3(x[1]),
    .I4(x[5]),
    .I5(x[7]),
    .O(_038_)
  );
LUT6  #(
    .INIT(64'hbcd399f6936c55ff)
  ) _091_ (
    .I0(x[3]),
    .I1(x[0]),
    .I2(x[2]),
    .I3(x[1]),
    .I4(x[5]),
    .I5(x[7]),
    .O(_039_)
  );
MUXF7  _092_ (
    .I0(_038_),
    .I1(_039_),
    .O(_036_),
    .S(x[4])
  );
LUT6  #(
    .INIT(64'h321348a51dd1dd33)
  ) _093_ (
    .I0(x[3]),
    .I1(x[0]),
    .I2(x[2]),
    .I3(x[1]),
    .I4(x[5]),
    .I5(x[7]),
    .O(_040_)
  );
LUT6  #(
    .INIT(64'h0bd0c3425695eb96)
  ) _094_ (
    .I0(x[3]),
    .I1(x[0]),
    .I2(x[2]),
    .I3(x[1]),
    .I4(x[5]),
    .I5(x[7]),
    .O(_041_)
  );
MUXF7  _095_ (
    .I0(_040_),
    .I1(_041_),
    .O(_037_),
    .S(x[4])
  );
MUXF8  _096_ (
    .I0(_036_),
    .I1(_037_),
    .O(y[6]),
    .S(x[6])
  );
LUT6  #(
    .INIT(64'h99600a55f03c0000)
  ) _097_ (
    .I0(x[0]),
    .I1(x[2]),
    .I2(x[1]),
    .I3(x[3]),
    .I4(x[4]),
    .I5(x[6]),
    .O(_044_)
  );
LUT6  #(
    .INIT(64'h3dcb71d4a3532f2f)
  ) _098_ (
    .I0(x[0]),
    .I1(x[2]),
    .I2(x[1]),
    .I3(x[3]),
    .I4(x[4]),
    .I5(x[6]),
    .O(_045_)
  );
MUXF7  _099_ (
    .I0(_044_),
    .I1(_045_),
    .O(_042_),
    .S(x[7])
  );
LUT6  #(
    .INIT(64'ha58196287bed7777)
  ) _100_ (
    .I0(x[0]),
    .I1(x[2]),
    .I2(x[1]),
    .I3(x[3]),
    .I4(x[4]),
    .I5(x[6]),
    .O(_046_)
  );
LUT6  #(
    .INIT(64'h4e723d7c39638ff8)
  ) _101_ (
    .I0(x[0]),
    .I1(x[2]),
    .I2(x[1]),
    .I3(x[3]),
    .I4(x[4]),
    .I5(x[6]),
    .O(_047_)
  );
MUXF7  _102_ (
    .I0(_046_),
    .I1(_047_),
    .O(_043_),
    .S(x[7])
  );
MUXF8  _103_ (
    .I0(_042_),
    .I1(_043_),
    .O(y[7]),
    .S(x[5])
  );
assign  { da[8], da[6], da[2], da[0] } = x[3:0];
assign  { db[8], db[6], db[2], db[0] } = x[7:4];
endmodule
